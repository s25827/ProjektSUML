��/      �xgboost.sklearn��XGBRegressor���)��}�(�n_estimators�N�	objective��reg:squarederror��	max_depth�N�
max_leaves�N�max_bin�N�grow_policy�N�learning_rate�N�	verbosity�N�booster�N�tree_method�N�gamma�N�min_child_weight�N�max_delta_step�N�	subsample�N�sampling_method�N�colsample_bytree�N�colsample_bylevel�N�colsample_bynode�N�	reg_alpha�N�
reg_lambda�N�scale_pos_weight�N�
base_score�N�missing�G�      �num_parallel_tree�N�random_state�N�n_jobs�N�monotone_constraints�N�interaction_constraints�N�importance_type�N�device�N�validate_parameters�N�enable_categorical���feature_types�N�feature_weights�N�max_cat_to_onehot�N�max_cat_threshold�N�multi_strategy�N�eval_metric�N�early_stopping_rounds�N�	callbacks�N�_Booster��xgboost.core��Booster���)��}��handle��builtins��	bytearray���B� {L       Config{L       learner{L       generic_param{L       deviceSL       cpuL       fail_on_invalid_gpu_idSL       0L       n_jobsSL       0L       nthreadSL       0L       random_stateSL       0L       seedSL       0L       seed_per_iterationSL       0L       validate_parametersSL       1}L       gradient_booster{L       gbtree_model_param{L       num_parallel_treeSL       1L       	num_treesSL       100}L       gbtree_train_param{L       process_typeSL       defaultL       tree_methodSL       autoL       updaterSL       grow_quantile_histmakerL       updater_seqSL       grow_quantile_histmaker}L       nameSL       gbtreeL       specified_updaterFL       tree_train_param{L       alphaSL       0L       	cache_optSL       1L       colsample_bylevelSL       1L       colsample_bynodeSL       1L       colsample_bytreeSL       1L       etaSL       0.300000012L       gammaSL       0L       grow_policySL       	depthwiseL       interaction_constraintsSL        L       lambdaSL       1L       learning_rateSL       0.300000012L       max_binSL       256L       max_cat_thresholdSL       64L       max_cat_to_onehotSL       4L       max_delta_stepSL       0L       	max_depthSL       6L       
max_leavesSL       0L       min_child_weightSL       1L       min_split_lossSL       0L       monotone_constraintsSL       ()L       refresh_leafSL       1L       	reg_alphaSL       0L       
reg_lambdaSL       1L       sampling_methodSL       uniformL       sketch_ratioSL       2L       sparse_thresholdSL       0.20000000000000001L       	subsampleSL       1}L       updater[#L       {L       hist_train_param{L       debug_synchronizeSL       0L       extmem_single_pageSL       0L       max_cached_hist_nodeSL       18446744073709551615}L       nameSL       grow_quantile_histmaker}}L       learner_model_param{L       
base_scoreSL       3.7122964E3L       boost_from_averageSL       1L       	num_classSL       0L       num_featureSL       24L       
num_targetSL       1}L       learner_train_param{L       boosterSL       gbtreeL       disable_default_eval_metricSL       0L       multi_strategySL       one_output_per_treeL       	objectiveSL       reg:squarederror}L       metrics[#L       {L       nameSL       rmse}L       	objective{L       nameSL       reg:squarederrorL       reg_loss_param{L       scale_pos_weightSL       1}}}L       version[#L       ii i}L       Model{L       learner{L       
attributes{}L       feature_names[#L       SL       citySL       typeSL       squareMetersSL       roomsSL       floorSL       
floorCountSL       	buildYearSL       centreDistanceSL       poiCountSL       schoolDistanceSL       clinicDistanceSL       postOfficeDistanceSL       kindergartenDistanceSL       restaurantDistanceSL       collegeDistanceSL       pharmacyDistanceSL       	ownershipSL       buildingMaterialSL       	conditionSL       hasParkingSpaceSL       
hasBalconySL       hasElevatorSL       hasSecuritySL       hasStorageRoomL       feature_types[#L       SL       cSL       cSL       floatSL       floatSL       floatSL       floatSL       floatSL       floatSL       floatSL       floatSL       floatSL       floatSL       floatSL       floatSL       floatSL       floatSL       cSL       cSL       cSL       cSL       cSL       cSL       cSL       cL       gradient_booster{L       model{L       gbtree_model_param{L       num_parallel_treeSL       1L       	num_treesSL       100}L       iteration_indptr[#L       ei iiiiiiiii	i
iiiiiiiiiiiiiiiiiiiiii i!i"i#i$i%i&i'i(i)i*i+i,i-i.i/i0i1i2i3i4i5i6i7i8i9i:i;i<i=i>i?i@iAiBiCiDiEiFiGiHiIiJiKiLiMiNiOiPiQiRiSiTiUiViWiXiYiZi[i\i]i^i_i`iaibicidL       	tree_info[#L       di i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i L       trees[#L       d{L       base_weights[$d#L       {�᠋�*��E_�"B�rEć�'E��D�i�m�#D�~�4�_Ľ�EmCfE�H�D�C��+��)C,E��D����z���A��НP�T��E�	SE8R�F�xE�m�D�=�E6�/C�o����F��!��D5zz��4�D�.eEQ��D<�Dąė��N}���C���ĭ%���č����yEa�SE��Ee�E{GoE�]EOVUE���E�D� �Db��E:�F��4�!�D>��1J��'��<C>1��|6�οC��D �ZBiFj¢3eC��sD#��D���D;��C�3�B���C�^�D-����ÚC$Ö�u�:]��;V��M�,Az)�C�;����ö<a��w�߄��ó���o ���)DSTD���DؓD�D�D�@�DbaD���E&�D��DpukD͍�DK��E�&C�uGD?w+B��C���C2'�DcN���BY�Ba�C��zB���s̱B�����+L       
categories[$l#L       B                               	   
                                        	   
                               	   
                            	   
                        
                             
            L       categories_nodes[$l#L       
                           #   <L       categories_segments[$L#L       
                             &       1       8       9       ?       @       AL       categories_sizes[$L#L       
                     
                                                 L       default_left[$U#L       {                                                                                                         L       idi L       left_children[$l#L       {               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c   e   g����   i   k   m   o   q����   s   u   w   y������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       {P���N�z�O�"No�NsHNߚ�M��KM6��L�xM��XM,3 M�=�M�@L���K���L9�8L���LYqPL��LK@L�V�L���L F`M��M%�0M�@M=s�Kї�Ka�KOEvJ��K�ǘK�-@L�TK�K�K�D�K% J�}�L� K~� K��`K��L&o\K�> L! K+�`K��L-n�L�O L�y�K�n�M-�     L�pL� L[�J��XJ�     J?�HKMLJ��@Jnݑ                                                                                                                                                                                                                                                L       parents[$l#L       {���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   5   5   6   6   7   7   8   8   9   9   ;   ;   <   <   =   =   >   >L       right_children[$l#L       {               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d   f   h����   j   l   n   p   r����   t   v   x   z������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       {B�        Bp     B�     B8  @�BH��@@  @@  @Z�HBճ3   @�@+�D�� D�  B        D�@ D�  B�  D�� B�  >���@S33B�  D�`    BG�D�` @ʏ\   ?���@�z�B�  D�  D�� Bl  B~B33D�� ?+�Bp  B�  ?ա�D�� D�� @�  EOVU?���=�hsD�� B�  >�  ��4D��    >Xb>H�9�<C>1��|6�οC��D �ZBiFj¢3eC��sD#��D���D;��C�3�B���C�^�D-����ÚC$Ö�u�:]��;V��M�,Az)�C�;����ö<a��w�߄��ó���o ���)DSTD���DؓD�D�D�@�DbaD���E&�D��DpukD͍�DK��E�&C�uGD?w+B��C���C2'�DcN���BY�Ba�C��zB���s̱B�����+L       split_indices[$l#L       {                                                                                             
                                                                               
                                                                                                                                                                                                                                                                         L       
split_type[$U#L       {                                                                                                                 L       sum_hessian[$d#L       {E�8 E�� D�� D�� Ev0 D/  C؀ Dʠ C�  E  D�` C�  C�  C�� C  De@ D0  B�  C�  D�� D.� D�` C�  C<  Cr  B�  C  Co  B0  B�  B�  C'  D;� C'  D@ BT  B,  B�  CC  D&� DC  C�  C�  D@ D`� CM  C  B�  B�  C  B�  B�  B  B�  B�  C/  B�  B,  ?�  A�  B,  BP  A�  C  B  C�� C�� C	  A�  C�  C}  A�  B  A�  A�  B  B`  B�  B�  C�  C�  C̀ C�� CY  C[  CF  B�  CK  C�  D� C�  A`  C?  Bl  B�  B(  A�  B�  @�  B�  B  A�  B�  B  B8  A�  Bd  @@  B|  C  B(  A`  BH  ?�  B(  A@  AP  A�  A�  @�  B<  A`  A�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       123L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       }@dOf���fE5ź�#6C���Et�Du�����+Đ��D�.��ô)ER��E���D���At���;pC�l�Ĭ���x]D�;�D(_C/���{ZE	�Et��E���E��
D��jE��C��ýgué�.C-׍�<�Oëf�Đ�7ĺsEč���8�"D��eE�B��Dn��D. ��[�"�B��	EX;QDס�E��EE'ɳE�@hDr/E�DE�e,DR��D�dD��E#ΚB�=D�`��	:�²���h�[�,�eCQ(:Ax�;Únc�J�z�vwB�3���ā�Ñmf�Ꝃ��G�ë��B��T�y�Z�%�!Dh C�)D�D��B�3�d.C/�C�lBRJC��ºĜB9�s^�w�B�)�����D-��D�׌C��~D&0�D�N�E��D>Dr��Dr.EzD��D�2E�DGܨC���CF�D:�Cf]C�SID7,DOuBc��;��C��B��"C� ��E��@��ڈB��XL       
categories[$l#L       Z                               	   
                               	   
                                     	   
                                  
                                           	   
                                  
                                           	   
             L       categories_nodes[$l#L                         
                  -   :   >L       categories_segments[$L#L                                    &       1       5       ?       B       H       I       J       K       L       YL       categories_sizes[$L#L                     
                            
                                                        L       default_left[$U#L       }                                                                                                      L       idiL       left_children[$l#L       }               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c   e   g����   i   k   m   o   q   s   u   w   y   {��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       }P {�N�\SN�ۼNlN��N*��Lܢ(Mu LP�`M�HL��M��M�Kҁ�K*y�L��XLw�@K\>�K�M�M
�pL��LD@�K�0L��M4�LI� L*�@K�shJ�#�K��I�vLƞK⭐K�$`LQtJ�� J�Y�K � J��K�y�L��@J��K�`L��K79nJ�P J�L��K�a�M/֠K�-�L0     K�k@K? J�аKpʠJ���J��PK ,J\7�I�g0I�M,                                                                                                                                                                                                                                                        L       parents[$l#L       }���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <   =   =   >   >L       right_children[$l#L       }               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d   f   h����   j   l   n   p   r   t   v   x   z   |��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       }B�  Bf           B�        B  @�   B�  @VffBճ3   BD  B@     D�� D�@    @�RD�@ ?�(�@�p�A`  D�@ D�` >�z�   >�(�   @@   @1G�B
ffD�� A�  BDp�D�` B�33>n��B��=B~B�     ?��D�  D�  D�� D�  >�
=Dr/=aG�A   D�� >���A�     B�  ?�7LB�     �h�[�,�eCQ(:Ax�;Únc�J�z�vwB�3���ā�Ñmf�Ꝃ��G�ë��B��T�y�Z�%�!Dh C�)D�D��B�3�d.C/�C�lBRJC��ºĜB9�s^�w�B�)�����D-��D�׌C��~D&0�D�N�E��D>Dr��Dr.EzD��D�2E�DGܨC���CF�D:�Cf]C�SID7,DOuBc��;��C��B��"C� ��E��@��ڈB��XL       split_indices[$l#L       }                                                                                                     	                                                
                                                                                                                                                                                                                                                                                                          L       
split_type[$U#L       }                                                                                                               L       sum_hessian[$d#L       }E�8 E�X D_  E�` D�� D� C�� EP� D�� D	@ D>� C�� B�  CY  B�  D�` D݀ D"  D]@ C�  Cs  C� C�� C  C�� B   B�  C-  B0  BD  B  D�@ C� D�� D� C[  Cր D  C�� C0  C  B�  C!  CC  C�  Cv  B�  B$  B�  Cg  B�  B  @   BT  AP  B�  B�  A�  A�  B  A0  A�  Ap  D+� C�  B�  C�  C�  Dk� C�  C�� B�  B�  C�  B�  D  @�  CQ  B�  A�  C  B�  B0  B(  B   B�  B�  B�  B�  C  B�  B�  B�  B<  A�  A�  A�  Bt  BP  CN  A�  B@  B@  @   B  @�  B@  A0  @   BX  B(  Bd  A�  A@  A�  Ap  ?�  A�  A   @�  @�  A�  @�  A   @�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       125L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       @���ùc�D̒-�F���>��E�C�#ö��C�%�Z��
lD�^�EX�DiֹB���*[�Ö��C����Ɯ��r'e�-�^�!�(E��D��)EBi�E��VD7m D���C�-�Ê*�����A7��ãf���D���3��Ò�CG��Ď"��b���a���@���A@�:���SoD'(Dں\E? $D���D��E'�E��8Dؙ
E���C��`D���C��%D���C�C�Bñ�pB��s�h���;Ã��G&�0��±�\�4�ZB�	C �_C���S��B`9)���BU'�C�n�U Wî�À��c�Ó]p�tӧâ{'�����RA�®H��>4��)�~%�¢�BO���%��Cf��C��DDn03D���D	V�C�W}A�LsB=�xC�3�D�6|D�DǨ3DmҵË�EDD��C�|sD� xB��vC���C��C�0�C���ϣmC�k�DI}C6��U�¹0'B���£��7;�B����6zL       
categories[$l#L       X                      	   
                                     	   
                               	   
                                           	   
                        
                         
                                     
                      
                      L       categories_nodes[$l#L                                  "   '   (   )   *   ,   :   ;   >L       categories_segments[$L#L                      
              $       2       9       @       A       B       C       D       J       K       R       S       T       UL       categories_sizes[$L#L              
                                                                                                                L       default_left[$U#L                                                                                                           L       idiL       left_children[$l#L                      	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c   e   g   i   k   m   o   q   s   u   w   y   {   }����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       O�}�M�\N�uDM[�YL*>�NA�L�~+LPM�L���K��@K�R@L��PM(7�K�D�Kլ�J\�@LNtDLWh"L�}J� J�`KU�JtrTL;��L�M��L���K��PKX��J�-J>?HJ�4�I�� K�N�K��L���J��Kzw�K�2I.� J���I�
 J� J��(J�� J�vI�ӀK�hL�K�i K�?L�� L^l�K�LI~@J��KvK`I�FJ�� J��J�B�I�l�Ie�d                                                                                                                                                                                                                                                                L       parents[$l#L       ���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <   =   =   >   >L       right_children[$l#L                      
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d   f   h   j   l   n   p   r   t   v   x   z   |   ~����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       B��=      BH��BDp�B�=q   @      D�  D�` @�D�@ B�Ǯ   @L(�A�  @�G�D�� @   B{   @T��      C  @   @�  @�  ?xbB�  A�  D�` D��    D�@ @@  BD  >��            ?CS�   @�  BH��?�Q�?.�A8��>���?:^5@�{>�u=��-D�� D�� ?�A�      ?��>��j   �h���;Ã��G&�0��±�\�4�ZB�	C �_C���S��B`9)���BU'�C�n�U Wî�À��c�Ó]p�tӧâ{'�����RA�®H��>4��)�~%�¢�BO���%��Cf��C��DDn03D���D	V�C�W}A�LsB=�xC�3�D�6|D�DǨ3DmҵË�EDD��C�|sD� xB��vC���C��C�0�C���ϣmC�k�DI}C6��U�¹0'B���£��7;�B����6zL       split_indices[$l#L                                                                                                       
                                             
                     	                              
                                                                                                                                                                                                                                                                       L       
split_type[$U#L                                                                                                                     L       sum_hessian[$d#L       E�8 E�� D�� Ez  D�  DG  D� E(� D�� D�@ D� C�  C�  Cq  C�� C�  EP D$� D � DB  C�  Cހ B�  B�  C�� C�  Bp  C-  B�  C1  B�  C_  Cg  D�� D� CՀ Cg  CÀ C|  CL  D  B�  C�� C:  C�� B�  @�  B|  B�  C�� B`  CR  B�  A   BP  B�  B�  A@  B`  B�  BL  B�  A�  B�  C  B�  B�  D  D�� Cр C  C�  B|  B�  B�  C�� Bx  C  B�  C6  A�  CD  C�  B�  B  B�  CE  B�  B�  B�  C2  B�  A`  @   @�  BL  A@  B(  A�  C�� A@  B   A�  B�  B�  B  A�  @   @�  @�  B@  B�  AP  A�  BT  A0  ?�  B  A�  B�  A�  A�  A�  B�  A�  A   AP  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       127L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       }@�R�NG�D���ß��C��aD���DX�E���F�D)&^����D��sE%4�DE��B->Ï!SAﻐ�Ã�"D��OC� ��5��C�aD��(DvCE`%bE��D��pD���C��ÜUFC.��C�:Lq�����/����O����D<�`D���C���D���B=2'ßv�B�C'D��D�i9��p�D45D��]Eq��C2�D�q�EcD0WDεXD�C�G1�d��C��t��,�DDJ�����Y��tC�!�C[�kB^�*®��A:a+���5npÀ�|�E��B�å�d]�0�~°��C�+�C$�mC��D-ŊC��#B�"C��*���ZC�5� Z����B��Q�;KeCr����uCz�D#{��i+DCW�BX�C�6C�+�Dy�\D�-D��X�r��C��Ci&�D��8DR-C�K}B��C�ǙB��D	��CAY����3Bnz���Y@���C�zI�f�gBN��C{xqB��aL       
categories[$l#L       s                               	   
                                     	   
                                        	   
                                  	   
                                            
                	   
                            	   
                               
                                  
                                   
            L       categories_nodes[$l#L                         
                     -   .   ;   >L       categories_segments[$L#L                                    )       5       6       7       8       9       ?       G       R       S       \       f       gL       categories_sizes[$L#L                                                                                                  	       
              L       default_left[$U#L       }                                                                                                         L       idiL       left_children[$l#L       }               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c   e   g   i   k   m   o   q   s����   u   w   y   {��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       }O�iM�� M�c$M�M�JMP��L�RLU<LI?�LE�XK�RLG� L��pKH/0J�WVJ�V�L'�K�G@K�q�Lz�L�2KK�Kk�tLgK�J`L�M�Lh>@K?�(J���J�b�J(�xJ�U@J��JK~!<K���K5� JzN�K�wK#\�K<L�K��(K���K�ԤKTJ��\J���KDn~L!$ J�x;K�)�L �@Le@J�Ll��K�z@J�[�J�G J��H    J��TJ��VH�B�I�-�                                                                                                                                                                                                                                                        L       parents[$l#L       }���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   ;   ;   <   <   =   =   >   >L       right_children[$l#L       }               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d   f   h   j   l   n   p   r   t����   v   x   z   |��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       }B�  Bp           B�     B      @�   @Z�H?2�      B�  @+�      D�@ D�@    A�  A@  ? Ĝ   B�  A�  @8�B�  ?�7D�� ?G�=D��D�� D�� @   ?}p�B  >B�\<�/>-V?�E�>\B|        >�B  B�  A   >?|�D�� D�� @�  D�` =��P@�C�G1   >���@�     �����Y��tC�!�C[�kB^�*®��A:a+���5npÀ�|�E��B�å�d]�0�~°��C�+�C$�mC��D-ŊC��#B�"C��*���ZC�5� Z����B��Q�;KeCr����uCz�D#{��i+DCW�BX�C�6C�+�Dy�\D�-D��X�r��C��Ci&�D��8DR-C�K}B��C�ǙB��D	��CAY����3Bnz���Y@���C�zI�f�gBN��C{xqB��aL       split_indices[$l#L       }                                                                                  	            
      
                                 
                                                                                                                                                                                                                                                                                                                           L       
split_type[$U#L       }                                                                                                             L       sum_hessian[$d#L       }E�8 E�X D_  E�� D�  D� C�� D�@ EJ� C�� D'@ C�  C�� CD  B�  D  D�� E
� D  B�  C�  C�  Cu  C'  C  B�  C*  Bp  C  B�  A�  D  B   C�� D`� D�` D.� C�� D� B�  BP  C�� B�  C  C�� C*  B�  C  Ap  B�  B(  B�  @�  B@  B�  A�  A�  C  @�  Bt  A�  A0  A�  C�  C�  A�  @�  B�  CO  C�� D� D�  B�  C  D
� B�  C�� C7  C�  A@  Bl  AP  B  B  C�  B|  A   @�  C  B�  C;  B�  B�  B�  A0  A�  C  @�  A   B   B�  B  A  A   B�  @�  @   B4  @@  B�  B  Ap  A�  @�  A�  B�  A`  A�  B,  A@  @�  @�  @�  A   A   L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       125L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       @����FZD����VE�C�DD�_�C��<����Ø�`D:�B�kID�8�D]*�D2�zB�G�Q>���ŋ�>Q�C�IDQ]��4T�C��2Do[aD��[Ci�%D�,rDM�$C��IB3�á\�C]Y~W�Ì����`ÁU�����Ô9�� |�Du&)C?�C��D���B&���x�#Dd3B�HB�&D�a�E�DE���m�D�u3D"��E#D/��DՆ�CwsD���C�S����C�����.@]�YB����xB���@����LA/���D�¯-�A�S�� Ѧ�ڷK��S��2����;�C(jCՇ�B
<A��C[ A�~'Cq�!C�T�D7�NBC/&�4��C�U­�J�'�CDkCQu7@�[Cn5�A=HC�WAؕ�D7�C�9�B��xC����jC;!+Cl1�Da%�C�UB�w�D;îA�p�C�c�B��tD8$C{��BjګCՖOB�,�D#�C?����_�¹fFAf��C��A�����8
�8�1L       
categories[$l#L       N                               	   
                                        	   
                                        	   
                                  
                             	   
                                   	   
                  L       categories_nodes[$l#L                                           =   >L       categories_segments[$L#L                                    *       +       3       4       5       6       7       =       >       LL       categories_sizes[$L#L                                                                                                  L       default_left[$U#L                                                                                                                    L       idiL       left_children[$l#L                      	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c   e   g   i   k   m   o   q   s   u   w   y   {   }����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       N��Ml�M#)�L���L~n�L�� Ku��K�9HLe�LA0K��LJ}�LO�zK%I�	GK��J�tKT�K��K̈́�LJ��J��K��K��|Ll�L�7LlJ��J��2Ik��I��.K��vKJ8JL�0J��J��K � J��pK}�1K�3�Kf�,K`4K�րJѷJo�PK��JL�K$��K(�Lq��K�K_�KG�0K4E�Ln J��I|�J��]J/ƄID��H�f`G��4I�:�                                                                                                                                                                                                                                                                L       parents[$l#L       ���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <   =   =   >   >L       right_children[$l#L                      
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d   f   h   j   l   n   p   r   t   v   x   z   |   ~����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       B�  Bx                    D�` D�  D�� @   D��       @�Q�D�     B4(�D�  A�     @a�>��yA@  C  >ɺ^@I�B�     >KƨD�` @@  @hQ�?��@@  B'
=A�  BX  ?BJ>�`BD�@ Ap  ?S��?�>49X>��?�@�  >vȴ>\(�A   >�\)>J��A�?S�@�  @�1>Z�>�M�>P�`      @]�YB����xB���@����LA/���D�¯-�A�S�� Ѧ�ڷK��S��2����;�C(jCՇ�B
<A��C[ A�~'Cq�!C�T�D7�NBC/&�4��C�U­�J�'�CDkCQu7@�[Cn5�A=HC�WAؕ�D7�C�9�B��xC����jC;!+Cl1�Da%�C�UB�w�D;îA�p�C�c�B��tD8$C{��BjګCՖOB�,�D#�C?����_�¹fFAf��C��A�����8
�8�1L       split_indices[$l#L                                                                                    
                                 
                  	         
                           	   	      
            	                                                                                                                                                                                                                                                                           L       
split_type[$U#L                                                                                                                         L       sum_hessian[$d#L       E�8 E�@ D'� E�� D�� C�  CE  D�` E^� D� D  C�  C  C   B  D�� D� E  D�� C�  C�  CЀ C?  Bh  C�  B�  B�  B�  B�  A�  A�  D� D@ C�  C1  D@ D�` D`� D  B8  C^  B�  C  C�� B�  B�  B�  A�  B  Cj  B  Bd  A@  B  B,  B�  A   B�  @�  @�  AP  @   A�  C�  C�� C� Bh  C  C�� C  A�  D  BT  D%  DK� D @ C�  D@ B,  A�  A�  C:  B  B�  B4  B�  A�  C4  B�  @�  B�  A�  B�  @�  B�  A   A  B  @�  CE  B  A�  A@  B0  AP  A   @�  A   A�  B  A   B  B  @�  @@  B�  @   @@  @@  @@  @   @�  A   ?�  ?�  @�  A   L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       127L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       @�f��8D$8��Q�AHwDgA�C^DK�hï�LB��X���D@�AD�%�C�7!��Û�|��lt�mt����wCVT[��˪�y���o��D0EݢE�0D�BC�O�DLq��[4�As�J�Fæ]��qS�9�Nµo\Ù_$����ñ�Cm�Ds��%�Cc��Ç�2C
b��︑C'�>D��C��^E:�C uD� OEN�HE�
DOu~A�EC�%(��D��$Ã��C��L��(\C8]�C�a�W�����Nª4B�V�����M®'t��?A2�`���B7�I�R�����Z3�S~Ap"^C ��A��CJ����w�B�.0´N$�|_?���CѨ��NC���1`�B����B�OC��C1m���s C�h�D��Ë]FC��#��]�D�8��TZD��PB�o�DLf�ÁºC��oB�
��C�oSB�`�£�C ��C�/_Cg������ �C �A���B����r��B������L       
categories[$l#L       k                               	   
                               	   
                            	   
                               	   
                                    
                                                           	   
                               	   
                               	                         
            L       categories_nodes[$l#L                         	   
            !   "   +   ,   2   3   <   =   >L       categories_segments[$L#L                                    #       .       /       0       1       7       8       <       A       D       J       W       X       Y       Z       _L       categories_sizes[$L#L                     	                                                                                                                       L       default_left[$U#L                                                                                                                L       idiL       left_children[$l#L                      	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c   e   g   i   k   m   o   q   s   u   w   y   {   }����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       N�PL�r4L�� K�ʨLV�L��HK� Ks��Js�K�(%K	��Lk'�L�K/I�JJZ KiP,JVJ�@K��J�jJd�J��(L/V�K�z�L��K��K�J�I���JW5JN:Is@JТ�J�L�I�dIH��I�� J�K���K-�JDIJ�+�J&�xI���J�D�JļCL��LK�K��K!��L�lKF��Ky��Kd� J~ԒJ�I7b.JS�I�"GAv�I�{I��L                                                                                                                                                                                                                                                                L       parents[$l#L       ���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <   =   =   >   >L       right_children[$l#L                      
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d   f   h   j   l   n   p   r   t   v   x   z   |   ~����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       B�  B@�         B�     @            D�� @VffB�  B�  ?fff@Vff   D�  BX  D�� D�� B�  @Q�? �D��    =��>&�yB�  >���   D�`       @�  @�  @�  A   @�  >���@@  @�      ?�?m�h?��\B  @�        @   >�+=�9X>�z�=�;d@   B�  >��         C�a�W�����Nª4B�V�����M®'t��?A2�`���B7�I�R�����Z3�S~Ap"^C ��A��CJ����w�B�.0´N$�|_?���CѨ��NC���1`�B����B�OC��C1m���s C�h�D��Ë]FC��#��]�D�8��TZD��PB�o�DLf�ÁºC��oB�
��C�oSB�`�£�C ��C�/_Cg������ �C �A���B����r��B������L       split_indices[$l#L                                                                                       
                  	                                                     
                     
      
                                                                                                                                                                                                                                                                                       L       
split_type[$U#L                                                                                                                   L       sum_hessian[$d#L       E�8 E�� D�� E[` E@ D/  C؀ EP D�  D�� D}� D� B�  C�� C  C�  D�  Ct  DG@ Dw� C׀ C�  D  D  A�  B   B�  Cu  B  BL  B�  B  Cހ DW@ D�� B�  C%  C=  D  DI� C9  C�� BX  CӀ A�  C�  B�  CF  C�  A�  @�  A�  A�  A�  B<  B�  C,  @�  A�  B@  @@  B`  B,  @�  B  CX  Ce  C�  D@ D-@ C׀ B   B  B�  B�  A�  C   C�� B�  D� C?  B4  C  C@  C9  B   A`  C�� C  A   Ap  A�  Cր B�  B4  B�  B�  C�  B  @�  AP  @@  @   A   @�  ?�  A�  @�  Ap  @�  B,  B  B  A�  C  @�  ?�  A   A�  A�  A�  @   ?�  A0  B4  A�  A�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       127L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       u@���[�UDA��y�C S�C�D���K��Zb%C\ګ�z��C�̩D�O�D���DRP�B�����]�6D2
C�{B�{���_�Îw�Í�C��E �D!��B�D�}�D,��E+��C%��9�2U���)�}6�
��D"�CA���D�GC3g-C�¬DN�sR�C��Ö��C8�-B�[���D��µ��D�^E_.ô�0DL�D����z�E;��	D�D&D�1�C�D�_A7kUB�2�*/XB��C���]*���=1C�|�vL�m¦E��÷�B�*CbWB�C�bN�ul�B��JC!�B	ą�	�Cv��A�����F-A�+�C�����C<Wp�����cW�B�,gB��0C�X�C���6F���'CRE^D�c�C�ڮC������C�hª��Ó�BB�OSCO�D)�CɛT���:Cf�>��u�C�D	��L       
categories[$l#L       9                       	   
                                           	   
                            
                                
                            	   
                L       categories_nodes[$l#L       
            	   
            /   8L       categories_segments[$L#L       
                                           !       "       ,       7       8L       categories_sizes[$L#L       
              
                                   
                     L       default_left[$U#L       u                                                                                                    L       idiL       left_children[$l#L       u               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K����   M   O   Q   S   U   W   Y����   [   ]   _   a   c   e����   g   i   k   m   o   q   s��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       uM��sL���LVV�KXK�<8K�tLK���K���J��pKԊ�J��[KxtKnn�L3R�L"�KD�TKT��J���H/UK���J�5�JJX�I�� Jp��KN�K!pJԏ�K'��K�vpK{��KV8KW,YJ�~nJ�(KR7�J:� Jo*�G�!�    K�)tK>J�TJ�j<J5� J���I�%H    I���J�mAK��I�LH�TJ���    J�+�JL`�J���Kc�K�.K���J��                                                                                                                                                                                                                                L       parents[$l#L       u���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   $   $   %   %   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   /   /   0   0   1   1   2   2   3   3   4   4   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <L       right_children[$l#L       u               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L����   N   P   R   T   V   X   Z����   \   ^   `   b   d   f����   h   j   l   n   p   r   t��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       uB�Ǯ@@           C  ?.{@
�HA�        =���@VffD�� D��    D�  D�` B@�@�Q�   D�@ A�  >j~�   >(��@_\)>%�T>j~�C  ?Hr�D�� @�  D�@ Bu�R@���B{B"��A���?z�D�� ?��B�  ?
��A  >bNC8�-   ?z�D�� >�+C  =�/ô�0@   C     =��
B�  @�  >k�C�D�_A7kUB�2�*/XB��C���]*���=1C�|�vL�m¦E��÷�B�*CbWB�C�bN�ul�B��JC!�B	ą�	�Cv��A�����F-A�+�C�����C<Wp�����cW�B�,gB��0C�X�C���6F���'CRE^D�c�C�ڮC������C�hª��Ó�BB�OSCO�D)�CɛT���:Cf�>��u�C�D	��L       split_indices[$l#L       u                                                                                         
                                     
                  	                
                                                                                                                                                                                                                                                               L       
split_type[$U#L       u                                                                                                           L       sum_hessian[$d#L       uE�8 E�h C�  E�( D�  C�� Cs  E60 D�@ D�@ D� Cf  B  B�  C  DJ@ E� D�` @�  D� D(  C�  B�  B  CA  Ap  A�  A�  B�  C  A   D  C�� D�� D/  D�  C�  @�  ?�  C�� Cq  C�  C@  C�  B�  B�  ?�  Ap  A�  C  B  @�  A0  ?�  A�  @�  A0  B�  @�  B�  A�  @�  @�  C�� CA  C�� A�  A@  D�@ D-� @�  D�  B$  C  C�  @   @�  C�� Bx  BT  C<  B   C�  C;  @�  B�  C�� B�  @�  A�  B�  @@  A@  A�  @�  B�  BL  @@  B  ?�  @@  @�  @�  AP  @�  @�  ?�  @�  @�  A   Bp  ?�  @@  B�  B  @�  Ap  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       117L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       w@�?����D	�¯�tB��C�NbDGF��%�>��Ar�pCY�[B���DftD��D�Bl�����®$�B��Bڠ��_���L5�C�$�C� �=rCͨqD�vQDv 1D���D��D�L�]òC���+���#\�� �S�K5�C]�T��<�C!������<��AZo�C}Mv��.�C*�;D!IA�V�D�1��]��BK�DA��C�E�MD93�â�TD�DGvÛ�`E�D�4�%Z�BWg�B�0$C�8��eA�7�fO��Z�@��@0Y1�ι(�,���B��N�7�VB�a�B��gB:<¯Q����� ��;�B<��>�<çtB�0G��6C���A��B���C%C�9cC�d�x(C�)A޶î8B	&�B�m8�&��C�R�Bh�B��}�ԶDc�=C�Z��d�C�8�y9B��]D(�Cv=WB�,�Crq6C���D<\C[K��� L       
categories[$l#L       !                                
                            	                            
                     L       categories_nodes[$l#L                                        *   3L       categories_segments[$L#L                                                                                             L       categories_sizes[$L#L                                                        
                                   L       default_left[$U#L       w                                                                                                     L       idiL       left_children[$l#L       w               	                                    !   #   %   '   )   +   -   /   1   3   5����   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c   e   g   i   k   m   o   q����   s   u����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       wM"L ZRK�~K���K��^K���K���KʄK3��J늴K�gcK1�MKBLK�bxK�V�J���J�� J|��K��JĊ�J�\J��K��8K�Z K=��J�?vK0�    K�K|K9��J�g�JC/�J�(KJߜ�J��xJE�TI���K�JO�J��bI�bJrDbJ�5nJ�RK�.KF��K3�tK1`wK*�zJ�@�K�{K|uJ��*J��0J��JCK��KC+    J<�H��p                                                                                                                                                                                                                                        L       parents[$l#L       w���                                                           	   	   
   
                                                                                                                                   !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   ;   ;   <   <L       right_children[$l#L       w               
                                     "   $   &   (   *   ,   .   0   2   4   6����   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d   f   h   j   l   n   p   r����   t   v����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       wB�Ǯ@@           B�  =�\)=t�A�  ?Y�>.{=�x�>�p�   D�@    >��         D��    A�  >�$�>cS�   >B�\Dv 1D�� A"�\C  BH��Ap  B   D�  D�@ >��D�� >�Z>$�/>t�B�     D�` @�  D�� >���@   @I��?��>�F   @ÅD�@ ?�ZB�  >C��>�=qÛ�`>�$�C  �%Z�BWg�B�0$C�8��eA�7�fO��Z�@��@0Y1�ι(�,���B��N�7�VB�a�B��gB:<¯Q����� ��;�B<��>�<çtB�0G��6C���A��B���C%C�9cC�d�x(C�)A޶î8B	&�B�m8�&��C�R�Bh�B��}�ԶDc�=C�Z��d�C�8�y9B��]D(�Cv=WB�,�Crq6C���D<\C[K��� L       split_indices[$l#L       w                                                   
                           	      
                               	                                       
                     	   
                                                                                                                                                                                                                                                  L       
split_type[$U#L       w                                                                                                           L       sum_hessian[$d#L       wE�8 E�h C�  E�( D�  C�� Cs  EI� D�� D�� D*@ C  B�  BT  C>  Ce  E;� D>@ D;@ C�� D$  B�  D� B�  B�  B�  B  @�  B@  C0  A`  C#  B�  C�� E� D� CZ  C�  CЀ C�  B�  Ca  C׀ A�  Bh  C�  C  BT  A�  A�  B\  B  B<  @�  A�  @�  B$  C,  @�  A0  @@  B�  B(  B|  @@  CG  C�  D�` D@  C  C�  B|  C  B  C�� C�  A�  B�  C�� B  BP  C<  B  C�� C  @   A�  BX  @�  C�  C  B�  A�  A   B,  Ap  @�  A`  @�  B  A�  Ap  A�  B  AP  @@  @@  @�  A�  @�  @@  Ap  A�  B�  B�  @�  @�  @   ?�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       119L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       {@m��#C���B�¡�QC�DB�;��|�B��T�$z��@�B��_C�HJD.l@���Å���#`����CF� ��>���Aɧ��aHD���:�C�cD��,CS��D�#�¿��C� a÷�LB���Af�B�dB�n}CɎ�B#SWC�������\F�A�����:@$��Ds�;�,CY4lC��D�|Cm�X���+C�	EDJ�E��C���~m�D]yD��K@��H�C�=D�2(Bd�N�(˨ BC>D"�c@�6�SB,�������BE�3� iuC���B�-C
����A�5�C8E������?wʉ�A�9��u�=�u���OWq�-�A��C�{�B�[T�%��3��yٙC��
D7r@����gC���O�CU*tC�KBGH�CЩC�w�C(47D7��X�C]s���5B���C� v����DsCzCc$��8C�`�-@��D!�<B�ɷ)L       
categories[$l#L       T                            	   
                                 
                                   	   
                                                        	   
                                           	   
                                        	   
             L       categories_nodes[$l#L                               '   ,   0   7   8   <L       categories_segments[$L#L                                                         #       $       )       7       E       F       SL       categories_sizes[$L#L                                                                                                  L       default_left[$U#L       {                                                                                                         L       idiL       left_children[$l#L       {               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [����   ]   _   a   c   e   g   i   k   m   o   q����   s   u   w   y������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       {L�r>K���K��XK>NyKe�K�v�KƾJV=(K��J�sJe�@K]�K]��JƑtJ�x�J �Jl>K5�K�:�Iǡ@J��J)�J�PKk�QKE|KJ��K8e�J!A�I�/�J��%KW'tI���J)��J:�I� �J�K�Jr�0KƵK��I�}^Id� J�xJ�@J��H��J�`    K,șK��K�]Kr�kK2��K�J@J]-0J:�IP�Iۥ�I�W`    JdD�J��<KKLJ�7�                                                                                                                                                                                                                                                L       parents[$l#L       {���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   ;   ;   <   <   =   =   >   >L       right_children[$l#L       {               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X   Z   \����   ^   `   b   d   f   h   j   l   n   p   r����   t   v   x   z������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       {B�        B,     D�@ >��A�  A�  B\)?�RD�  A�  ?�G�>�ff@�p�@�  D�� D�� >�5?   @�  AP  >�ȴ   B�  >��>q��   ?M�?��   A0  B33?�ȴ>�t�>w��D�` ?%�   >�`B@a�D�� @      @�CY4lB̊=   >�jC  @Z�H>C�>%>["�      =�Q�@�D�    D�  D�` �(˨ BC>D"�c@�6�SB,�������BE�3� iuC���B�-C
����A�5�C8E������?wʉ�A�9��u�=�u���OWq�-�A��C�{�B�[T�%��3��yٙC��
D7r@����gC���O�CU*tC�KBGH�CЩC�w�C(47D7��X�C]s���5B���C� v����DsCzCc$��8C�`�-@��D!�<B�ɷ)L       split_indices[$l#L       {                                                                                   
                            
                
                                       
   	                                                                                                                                                                                                                                                                             L       
split_type[$U#L       {                                                                                                              L       sum_hessian[$d#L       {E�8 E�� DZ� E
@ Ey� D@ C�  D@� D�@ EP D�` C  C� A�  Cl  B�  D-� D-  D;� D� D�� C   D�` B(  B�  C�  A�  AP  A  C/  Bt  Bh  A�  C�� Cv  D  Bp  C�� C�� C�� C7  D�@ Cƀ B�  @   D�  @   B  @�  BX  BX  C�� B�  A  A   @�  @�  A   ?�  B�  BP  A0  BH  A�  B  @�  A@  C�  C  B�  C  B�  D� A   BH  BH  C�� C  Cl  C�  B�  A�  C&  DS  D� CH  CE  @�  B�  ?�  ?�  D�� Cm  A�  Ap  @�  @   B<  @�  B4  A  CM  C  A  B�  @   @�  @   @�  @�  ?�  @�  @@  @@  @�  @@  B�  A�  A�  @�  @�  A�  A�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       123L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       o@W����wC��3�_�jB��C��'��+|¼���i@�mC �BD `�C2���b%&D?l��ЖPB��a¸�]A���?��B���C���@w@Cl5D[IUC�m��
�Y�C��*B�n�C�k��I��%�ø�C$����BS���]B�+&CԍR�a�1B�RC��Cٞ�}�Ú6LBc��B	p1D�ˆD��yCb\�DH�SBq��V��Abf�C��Q�Bp����V����@�kC	�$�D����a4A!#�B���B^���uB�F��IZ�?f���Q{B��{@����ɓ?D0���P.���x�A����
�C���uM�CQb�B���µ\BR_�Cv��
�@�[mB����(�C�DL9zB�R��\��C��C�p��]#�C��?�����]�C��8�-h�����B�zzA�k-�>2�(m�L       
categories[$l#L       @                            	   
                         	   
                                                     	   
                                  	   
                              
                  	L       categories_nodes[$l#L             
               !   #   &   *   7L       categories_segments[$L#L                                                                       '       2       ;L       categories_sizes[$L#L                     	                                                        	       L       default_left[$U#L       o                                                                                                L       idi	L       left_children[$l#L       o               	                                    !   #   %   '   )   +   -   /   1   3   5   7����   9����   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c   e   g   i   k   m������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       oL6}KP�K{'xJ�tK�"K�\�Jk��J�ݸJ�s�J�HAK��K��\Kt݅J�Iq�8J0T�I���I��J�BmJ��Jߍ�KO�lJ^ݚK7f�K�>�K���J�BI��    G
    J#�mJ9`G�%HI�z�I�ݸJ��Jb@J�D�K��Jgs�J���K#<�J�UXJ�e�J<�J��Kn��Ke�WK�
�KZ, KH�lJ�|rJ�9dI�JN,GǛ�                                                                                                                                                                                                                        L       parents[$l#L       o���                                                           	   	   
   
                                                                                                                             !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8L       right_children[$l#L       o               
                                     "   $   &   (   *   ,   .   0   2   4   6   8����   :����   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d   f   h   j   l   n������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       oB�ǮBK��   @�  D�@ =��?��RB�  B  A�     D�� B  ?�ƨ      A�     D�� D�` A@  @��
>49X?ƨ@�  @�  >^5??���C��*   C�k�D�� =o   D�@    =���=\   B�  @���@j�H   @@  @   >�G�B�  @�  @�=��-=#�
>�{A�  >p��D��    @�Bp����V����@�kC	�$�D����a4A!#�B���B^���uB�F��IZ�?f���Q{B��{@����ɓ?D0���P.���x�A����
�C���uM�CQb�B���µ\BR_�Cv��
�@�[mB����(�C�DL9zB�R��\��C��C�p��]#�C��?�����]�C��8�-h�����B�zzA�k-�>2�(m�L       split_indices[$l#L       o                                            	                              
            
                                                            
                                                                                                                                                                                                                                                          L       
split_type[$U#L       o                                                                                                    L       sum_hessian[$d#L       oE�8 E�h C�  Ez  E � C�  B�  D�  E � E � C�� C7  CG  B�  @�  D�  B�  D.@ D�  D�@ Dx� C�� CZ  B�  B�  C.  A�  B�  ?�  @   @@  D!� D�  @�  B�  D  B�  DN  D@ A�  D�  D]� B�  C>  B�  A�  C;  B`  A@  B�  A�  B`  B�  A�  A  B�  A   ?�  ?�  C�  C�� A   D�  @�  ?�  B0  B  A�  D� A�  Bt  C
  D+� C3  C�  Ap  @@  Dz� B8  D+  CJ  B�  A�  Bd  C  B$  Bx  @�  A�  C)  A�  A�  B   @@  A  A   B�  A   A�  B,  AP  B�  @�  A`  @   @�  @�  B�  B  @@  @�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       111L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       q@2���
�B�MZ��@�|�C0A��y�C�/-���'�թB�E�C#�pD�8rAJcP���q��J�)lL���P�»0A��b��لB�j�Ch*<A���D�t�B�u��d<D���1c1CNZ:AD-�:D-4����J��m��Y�*��C'�����B��[�B�R��]�wC	�+�HC��?���5�k��B�x�B~4D��t�Ш{C ��zC��D[S"È�@^*�MAo����Z_H�@�\���·ÕC�����&��Bb�@K���T��ÆIw\�&�� �uBw�U�BSKB�l��&~B���?�������B ��B�����,#B�3�A�� B�����p�[W�BrT�C(:�CPP�����~Az��Q�wBU��C]_�Dq�,�����Ag1C	�%C�t��?�@H&g�)4����äHJL       
categories[$l#L       +                          
                          	                         
                            	   
                               L       categories_nodes[$l#L                            %   *   .   4   9   :L       categories_segments[$L#L                                    	                     $       %       &       '       (       *L       categories_sizes[$L#L                                   	                                                        L       default_left[$U#L       q                                                                                             L       idi
L       left_children[$l#L       q               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;����   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c����   e��������   g   i   k   m����   o����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       qK�9�J��K#��J@��J�¾K?��JppAJU�6J9G�J�l�J��KupJ�,`Jf�oJ�F�JD�xJ7�I�ڬJL�TJ�tIJ�JIg�JӣK1
�KM�I�X I���J��JM�)I)`    Jo$Jb-I�PI�&�Im��I��SJQI�DI��J@�,J�3�I��mJ!�I���J��&H�|KQd�J�|�J�3K/5    H��         JL��JzNJAhH��q    IA
(                                                                                                                                                                                                                L       parents[$l#L       q���                                                           	   	   
   
                                                                                                                                   !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   4   4   7   7   8   8   9   9   :   :   <   <L       right_children[$l#L       q               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <����   >   @   B   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d����   f��������   h   j   l   n����   p����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       qB�  A�        D�� A�  A&�\A��   >'�>�+>_;d?��D�� @@  D�� AP  >���@   D�    >�P      >ix�D�` >�7LB�  @��R>I�CNZ>���>��@H��@@  ?��7@X     @@  @�  >���D�     >�bN>��!Bh     ??}=�;d>��D�  B~4   �Ш{C �=�o?%`B      ^*D�` ����Z_H�@�\���·ÕC�����&��Bb�@K���T��ÆIw\�&�� �uBw�U�BSKB�l��&~B���?�������B ��B�����,#B�3�A�� B�����p�[W�BrT�C(:�CPP�����~Az��Q�wBU��C]_�Dq�,�����Ag1C	�%C�t��?�@H&g�)4����äHJL       split_indices[$l#L       q                                                                                                                                                     
                                                                                                                                                                                                                                                             L       
split_type[$U#L       q                                                                                                     L       sum_hessian[$d#L       qE�8 E�� D�� E)� E1� D�  C�  D�� D,� D�@ D}  D@ A@  C� Ap  D�  CG  Cڀ C~  D[� Do  C  DW� D,  C�� A   @�  C�  A0  AP  @   DS� Dt@ CD  @@  CZ  C[  A�  Cg  Bp  DL� C�  C�  B0  B�  D?@ B�  D� C  B�  Cq  ?�  @�  @   @   C�� C  A   @@  @@  A   C�� C�  BT  Dg  B�  B�  @   ?�  CL  A`  C7  B  A0  A@  CO  A�  Bh  @   A�  DF  C*  C�  C̀ BL  B   A@  B�  A   D%@ B�  A�  B�  C�  C  A�  B�  B,  BD  Ap  Cb  @   @�  B�  Ck  B�  A�  @�  @   @   ?�  @�  @�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       113L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       e@ ���(��C$���]-~C�F�C�G�B���@���dw�D7|�CWWeCb0D���B��-D8����BwKA�r���D9�B���D��C�D�/��IHCz�-�p��AOd�D�3��W�R�NB����h�Ä�B��):���hC��KDk��C}irÊ��Cz�� �C�-�D�}NA���� ��:Q�C�o����B� �
iC{�}CRkE�|A���˝�� µ�QA��D��A�%�x����yB�
B<�b����>X�����/�l�<8�B�����(�C���B��7B�����>���P�?dwM�C�O�f$�A�ק�:u�B���B&@C����5�CG�1C'���7V�o w�)J�V��B��A���)B� ��ǦgD7E9C2�]L       
categories[$l#L       4                            	   
                            
                                      	   
                                                          	   
   L       categories_nodes[$l#L             
            "   $   )   +   0   5L       categories_segments[$L#L                                                         $       '       (       )       3L       categories_sizes[$L#L                     
                                                        
       L       default_left[$U#L       e                                                                                      L       idiL       left_children[$l#L       e               	            ����                        !   #   %   '����   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U��������   W   Y   [   ]   _����   a   c����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       eK\i�J��pJ�4J�2�K�*K8�'J�o�J�xI��L    J��J���Jݐ�KKO��J�{�J���I��I�ˀI�pJd�-    J�JĨH2�KL+�K5UhI�X�J�"$Jk��I�{�K���J�k�I��.I�I�ڰIQ�|H3�I@��JRI�0�J���I"��G�VIڊ         J�IK1�>J1BlK5Y�IO�    G�&2Ip�                                                                                                                                                                                        L       parents[$l#L       e���                                                           
   
                                                                                                                                   !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   /   /   0   0   1   1   2   2   3   3   5   5   6   6L       right_children[$l#L       e               
            ����                         "   $   &   (����   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V��������   X   Z   \   ^   `����   b   d����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       eB�ǮA@  =�S�   =�hsD�� D�� @@  =�\)D7|�   B�     ?WK�?@  A"�\?tz�>"��   BH��B  D��@�{=<j   >\)>]/@�@   ?h��D�� ?r�!B�  >��#   =ȴ9   A`  >'�@��
@@     @�     ?���A���� �>���   >���?�  ?��C{�}   @�  A���˝�� µ�QA��D��A�%�x����yB�
B<�b����>X�����/�l�<8�B�����(�C���B��7B�����>���P�?dwM�C�O�f$�A�ק�:u�B���B&@C����5�CG�1C'���7V�o w�)J�V��B��A���)B� ��ǦgD7E9C2�]L       split_indices[$l#L       e         	       
                                          
                            	                                                                                                                                                                                                                                                                                   L       
split_type[$U#L       e                                                                                          L       sum_hessian[$d#L       eE�8 E�h C�  E�  B�  B�  C�  E�� D�  ?�  B�  BP  A�  C�  A�  ED@ D�  C�  D�  A`  Bh  @   BH  Ap  @@  CB  C`  A0  @�  E<p B�  D,@ D� A�  C�  D�� A   @�  A  B  A�  B0  @�  @   AP  ?�  @   BL  C  B   C@  A   ?�  @   @�  C�  E*� BH  B�  D*� @�  D  B�  A�  @   B�  CP  C  D�� @�  @�  @�  ?�  @�  @@  B  @�  AP  @�  A�  A�  @�  ?�  ?�  ?�  ?�  A@  B0  @�  B�  B   A�  A  A�  C.  @�  @@  ?�  ?�  @�  ?�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       101L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       i?�_���CA�e�&}�A��p�C%Cp�LC
��@�O�!��B`����D< �CN�%D��zÄ	�C�7��/PÃg��@� �BL~C���C��6��C�*eB�.�C���A�dhDk�C�'Cm� ��uFBf��C���IM�BՄ�æVJC�#×eA���BG�4A`B덜���D�=BN�eB�6³� à���ы��5��C9_�B�F�C���Ãg�C�����[�B=�h+�f5���o%B��jC���B�<�¤���\6�BQ�q�6[G�Ltg�"$��N[Cl�z�f:��;E��/'�Cڐ�@�#_BǢT��%���uA��=B���0A]�{��i�C^���k#Bʨ��@��A���B���-5���>Z�3 B��A� �HCDP�C@��A}0Z�Vs�A�1�CT��J�7L       
categories[$l#L                                          	   
                                               	   
         L       categories_nodes[$l#L                   "   4L       categories_segments[$L#L                                           L       categories_sizes[$L#L                                          L       default_left[$U#L       i                                                                                                   L       idiL       left_children[$l#L       i               	                                    !   #   %   '   )   +   -   /   1����   3   5   7��������   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W����   Y   [   ]����   _   a   c   e   g������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       iK	�J�eJ��JbsJ�n�J�|�K��J���J-�J��K2�J}�RJxJ�ϜG�S�I��sJxb�J2�
JAx>K��J�"K�K3|H��J�,    G<�zJ��2J�l�        HG��I��I�P@J���J+�XJ�-]Je��I��%J�l�J��.J�7�J�L�K'b�K c�K�J8�    GM0KI�7I��    D ��K�VJ�J���Ke\                                                                                                                                                                                                L       parents[$l#L       i���                                                           	   	   
   
                                                                                                                       !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   0   0   1   1   2   2   4   4   5   5   6   6   7   7   8   8L       right_children[$l#L       i               
                                     "   $   &   (   *   ,   .   0   2����   4   6   8��������   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X����   Z   \   ^����   `   b   d   f   h������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       iB�     ?�G�D�  >�C  B�  ?#�
B�  >�"�BP  >O�@�  >�   >P�`BX  @�  @BM�D�` >��P>� �>Y�   D�� C�*eD�� D�� >dZDk�C�'B  >��>s�F   =,1@�  B̊=>fffB�  Bճ3B�  >��
B�  D�@ ?&ff=���B�6B�  B�  B�  �5��   >��y@�z�A@  >\��[�B=�h+�f5���o%B��jC���B�<�¤���\6�BQ�q�6[G�Ltg�"$��N[Cl�z�f:��;E��/'�Cڐ�@�#_BǢT��%���uA��=B���0A]�{��i�C^���k#Bʨ��@��A���B���-5���>Z�3 B��A� �HCDP�C@��A}0Z�Vs�A�1�CT��J�7L       split_indices[$l#L       i                              
      	             	                                                       	   	                                                                                                                                                                                                                                                                        L       
split_type[$U#L       i                                                                                                    L       sum_hessian[$d#L       iE�8 E�� Ck  EC` Eh` A�  CR  B�  E<� D�� E � A�  @�  CN  @�  A�  B�  E8� Bp  C�� DM  E  C)  A   AP  ?�  @@  B�  B�  @@  ?�  @�  A�  B8  B  E1  B�  B\  @�  C1  C  D%� C  DZ  D�  B�  B�  @�  @@  A   @@  ?�  @   B4  B�  B   B4  ?�  @�  @�  A`  A�  A�  AP  A�  BX  E-� B�  A   A�  B  @   @@  C  B0  C  @   D  Bh  B(  B�  D(� CE  D  D{  A�  B�  Bx  A�  @   ?�  @@  @�  ?�  @   ?�  ?�  A�  A�  Bd  A�  A�  A�  A�  A�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       105L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       _?��B�M���9B+�D�H����+�C�EC���B���dX[B85��vT«�AD��B���B��Dr�7B8FB�������vk"����CdA�%9��]Bo��D4��Cq���C����e�iD�IDB��BG�}�)I�.�Cf���^ġs��ԥ�B46B0p�C�w�B�c����AUV\B<[t�źUDG�@�&gCB	B��Eª�HB���C��TBa�%�L�B.�"B#y6C���@7�pB����z+���9�
6���1-C-���XW�����K����A��#���2��@�BL�C<]�����B�}��'�A����Y����2�~��Ay#+��A�@�x��@C}.B�j�MBX*B�@�ٚL       
categories[$l#L       H                               	   
                                               	   
                                         
                            
                               
                         	   
             L       categories_nodes[$l#L                          +   ,   -   0   1   4L       categories_segments[$L#L                                                          ,       3       ;       <       GL       categories_sizes[$L#L                                                                                    L       default_left[$U#L       _                                                                              L       idiL       left_children[$l#L       _               	               ����                     !   #����   %   '   )   +   -   /   1   3   5   7   9   ;����   =   ?   A   C����   E   G   I   K   M   O   Q   S   U����   W   Y��������   [����   ]����������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       _J�oeJ�܄J@c�J˖?I���J!%I�K^Ku[�J�[BH�Ѡ    JQP)I���Ih"�IM�K�PKtnrJ���J!]-    I: I���I��6I��CI�D`G~�H�2PHz,LH�G�J��lJ��EJ�1*    J�FI��J��Jj    H` J�J(IN�JQ��I�j^I���I���I�B�    E��hG4�         F��    E�"�                                                                                                                                                                L       parents[$l#L       _���                                                           	   	                                                                                                                           !   !   "   "   #   #   $   $   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   0   0   1   1   4   4   6   6L       right_children[$l#L       _               
               ����                      "   $����   &   (   *   ,   .   0   2   4   6   8   :   <����   >   @   B   D����   F   H   J   L   N   P   R   T   V����   X   Z��������   \����   ^����������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       _   B�  A@  D� ?p��A   >A�7?S�A"�\=oB85�A     >��#   >�  B�  ?K�>�G����B8Q�@�  B6  ?<�A@     B�  D��    D�� D�` @@  DB��D�  B4(�B�  Bt  ��^D�� @   B�  =��`?@A�         B�  B<[t      @�&gCB	   ª�HB"��C��TBa�%�L�B.�"B#y6C���@7�pB����z+���9�
6���1-C-���XW�����K����A��#���2��@�BL�C<]�����B�}��'�A����Y����2�~��Ay#+��A�@�x��@C}.B�j�MBX*B�@�ٚL       split_indices[$l#L       _                         
                   
                                                                                                                                                                                                                                                                                                         L       
split_type[$U#L       _                                                                                    L       sum_hessian[$d#L       _E�8 E)0 E�� E(� A   E�� A�  B�  E!� A  ?�  EmP D� A@  A�  B�  A�  E  C=  ?�  A   Ei� B`  C  C̀ @@  A  A  @�  B  B<  A�  @�  E@ A@  C,  A�  @�  @�  EQ` CÀ A�  A�  B�  B�  C�� B�  ?�  @   A   ?�  @@  @�  @�  @@  A  A�  A�  A�  A@  A  D�  DZ� @�  A   C  A�  A  A   ?�  @@  C̀ E7� C�  AP  @@  A�  A�  A0  A�  B  A�  B0  C2  C  B�  @�  ?�  ?�  @�  ?�  ?�  @�  @   ?�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       95L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       a?��п�
'Cy���w{Al�$C�y��r��ŋw��Rp�OwuB�G$��#CC�Á��+B����7D��qz���t���N��@`Qo���C"��Ax�t��WDj�C�V]C�R�,�@����l8���2:���@���³�n� �p���Û�.C΁A���&�Y���D ���'��Cl1T�IZ
�BD�mm�l��B�ƩDW<6�?-�C/�B�����-��"�1¼�J�?i�B��Br���q/=��93@�I\�a�A��B�c��l�M�`��@�vU�Y.�J�Ci���Zꁾ�~B2�C1�+��
�!����C�'��%���	�}B���B���Cǒ>C�+�C��Ac���Bl}YÄ�B��C���Î	���V Cb��bR�L       
categories[$l#L                                            	   
                                   L       categories_nodes[$l#L                         0   3L       categories_segments[$L#L                                                         L       categories_sizes[$L#L                                                        L       default_left[$U#L       a                                                                                    L       idiL       left_children[$l#L       a               	                        ����            !   #   %   '   )   +����   -   /   1����   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S��������   U   W   Y   [   ]   _��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       aJ��JQ�kJ�I�Y�Jz��J��&K8}ItwhI���JAC�J�n�HΎPJ���    JJ�IpM�I-�VI�wI��J��J?.{J!"�J�Yh    G�6`Jdt�J��t    J+ÒI��I#�I2��IN�I��AI�t�I���It�0J,J+Jb��J��sI���J��J؃J�Vd        I���H�OJ?}�I��I!��I�D�                                                                                                                                                                                L       parents[$l#L       a���                                                           	   	   
   
                                                                                                                       !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   /   /   0   0   1   1   2   2   3   3   4   4L       right_children[$l#L       a               
                        ����             "   $   &   (   *   ,����   .   0   2����   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T��������   V   X   Z   \   ^   `��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       aC  B,  ?2-A��HD�@ =�C  >��#@��=,1A@     @�  ��+A   =�Q�D�� ?�^B  ?�V@�  B�  >��Ax�tD��    >�ƨC�R         D�� >.{=�
=?4�j=oD�� =�`B?��B�=q=���=<jD�� >�|�?9�#�IZ
�BA      >�J?
~�   D�@ B�����-��"�1¼�J�?i�B��Br���q/=��93@�I\�a�A��B�c��l�M�`��@�vU�Y.�J�Ci���Zꁾ�~B2�C1�+��
�!����C�'��%���	�}B���B���Cǒ>C�+�C��Ac���Bl}YÄ�B��C���Î	���V Cb��bR�L       split_indices[$l#L       a                  
      
                                      
                                                          	   
                  	                     
                                                                                                                                                                                      L       
split_type[$U#L       a                                                                                          L       sum_hessian[$d#L       aE�8 E�� B�  E� E�� Bp  A�  C�� EP E^` Dn  @�  BX  @   Ap  B�  CW  D�  C� B�  EY� C�  C�  ?�  @�  Ap  B  @@  A@  A�  B�  C"  BT  D�� Cl  C�� C  Bx  A   ES` B�  C� @�  B�  C�  @�  ?�  AP  @   A�  A   @�  A   @�  A`  B  B$  C  @�  @�  B@  Cx  D�� CS  A�  @�  C�� B�  A�  A   BP  @�  @�  ED  Cv  @�  B�  @�  C�  @@  @   B�  A�  C�� @@  A  @�  ?�  ?�  A�  @   @@  @�  @@  ?�  @�  @�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       97L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       W?]�BH�����B8r�D��]�>�hB�
A�J�C{��D5B���/��w�@Cf�R BQB��B���D{��T��C�g�����pBC>�D;���!ZD  ����B)V���çYPBZ��C�%�ETC�% �uĢ���C���å�Pîq�C���J�B��PC�v-B ðC`�WD��5¡_�+�&Dp�E¤E+�<â�|¹\�AvTA�Y���z��SGB�������(@V�P *@%�<��2mC<���@~ú���Z�B��;A�UCz@Q�X}�´�!CZ�����B�@��E9\CYNC�l�B��4�6�vB��Ö�RB�w�C�DM��| L       
categories[$l#L       $                                      	   
                                                              	   
         L       categories_nodes[$l#L       	                   #   '   (   +L       categories_segments[$L#L       	                                                                L       categories_sizes[$L#L       	                                                               L       default_left[$U#L       W                                                                        L       idiL       left_children[$l#L       W               	            ��������                        !   #   %   '   )   +   -   /   1   3   5   7����   9������������   ;   =   ?   A   C   E   G����   I   K   M   O   Q   S   U����������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       WJ6�J�
�J?�5JMovI�E\JTQCJ���JN�GJ�'�        J_GJ�=J�Q�J�'�J9RI��J��Jb�J�oKA��J���Iz��J:,;J�äJ.�2J[�_I���J9B1H�K�    I�            J)RrJ��K/�J���J�P�J%��H���    J��J�e�J	�HI��xJ�J:�lI�{�                                                                                                                                                    L       parents[$l#L       W���                                                                                                                                                                                   #   #   $   $   %   %   &   &   '   '   (   (   )   )   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1L       right_children[$l#L       W               
            ��������                         "   $   &   (   *   ,   .   0   2   4   6   8����   :������������   <   >   @   B   D   F   H����   J   L   N   P   R   T   V����������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       W   A�  B�        @�  @�  B�  @�  D5B��B�=q?MO�@�  >��j=49X   >��=��   @�  >gl�AP  >q��C  >��y?bNBx  =L��>�ZçYP>�I�C�%�ETC�%    >I�D�� A`        D�` B��P   D�� ?�{=���?:�HC  B�  ¤E+�<â�|¹\�AvTA�Y���z��SGB�������(@V�P *@%�<��2mC<���@~ú���Z�B��;A�UCz@Q�X}�´�!CZ�����B�@��E9\CYNC�l�B��4�6�vB��Ö�RB�w�C�DM��| L       split_indices[$l#L       W                                                   
                                           
       
                                                     
                                                                                                                                                          L       
split_type[$U#L       W                                                                              L       sum_hessian[$d#L       WE�8 D�� E�� D�� @   E�H CH  Dr� B�  ?�  ?�  E�` Bt  B�  B�  Dp� A   Bx  A0  E�( C  B  A�  B�  A�  B�  A  A0  Dn  @�  @@  Bt  ?�  @   A  Da@ E�  B�  B  A�  A�  A�  ?�  A�  B�  A   @�  Bp  A   @�  @@  A  @   A�  Dh@ @@  @   B  A�  D^� A   D�@ E_` B   Bd  B  @�  AP  A   A  @�  A�  @�  A�  A   B  B   @�  @�  @�  @   BT  @�  @�  @   @�  ?�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       87L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       s?D&�A>|��.@/]B���B��o�����ŵB�-B� |��3=B�D:N¼k���J2B�'a�_`Cػ_Bz��C���B��A�y�B�BB�o4�6t£q�Dh+@@�X��#���7C.Y�B��cD2B��\�4�&��D���B��B҉KcDNl�C.B=��C����J����F��.�Cw�PC,���'�~��J�ÇJQDz-2B�����NB����rS?k��a��xK����C��B@\#��q{B���C�!@$rT�ѳ���o群�C���A
[�OB���BT�4��.�A�Lq��PC�Ԯ��]�B�?VB�Z?;f��6C�lCC%Y�D'W�AI��G�1C���ZL5A�JEC1��B�WA�ir����°�C��B����0��BI�$A﯇�	�.��y�E��(�B��L��
B�f���Q��B�� Bg��C��L       
categories[$l#L       V                   
                                           	   
                                        	   
                                                             
                                      	   
                                            	   
             L       categories_nodes[$l#L                         !   $   %   ,   -   0   3   ;L       categories_segments[$L#L                      
              &       *       +       ,       -       8       9       F       G       UL       categories_sizes[$L#L              
                                                                                    L       default_left[$U#L       s                                                                                                     L       idiL       left_children[$l#L       s               	                                    !   #   %   '   )   +   -   /   1����   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _��������   a����   c   e   g   i   k   m   o   q������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       sJ"(HJ4$�I�J<�xJ�]*JW	�I���J=��J/r�J���JF8J�I��`J=YCI��6Jv�aJ)͜J��4J�J���J��JnJ#�I�;wH�s(    G���I���JS��JSJI��J,}�J+,�I��J1�I��8I�_hJ��I��bJS��I�P�JN�5J��I�+�I�� Jr.I�DIq�Hx�        H'�@    IsľI���Jn�DJ(5�I��)IU��Ib��I��V                                                                                                                                                                                                                        L       parents[$l#L       s���                                                           	   	   
   
                                                                                                                                   !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   3   3   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <L       right_children[$l#L       s               
                                     "   $   &   (   *   ,   .   0   2����   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `��������   b����   d   f   h   j   l   n   p   r������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       s>��h?M�=�t�D�� @2�A�  ?�D�  =��?�T>-V?|�B
ff   A/\)?�o=]/   ?U�   @�@�1?��      £q�A   D�� A�  A��@�  @@  >E��   >o��B�33      >�V=49X>>v�D�` @   <���      @�1>�{   ��J�ÇJQ   B��A   @�ƨB[��>�x�A
=?1&�   B\33B@\#��q{B���C�!@$rT�ѳ���o群�C���A
[�OB���BT�4��.�A�Lq��PC�Ԯ��]�B�?VB�Z?;f��6C�lCC%Y�D'W�AI��G�1C���ZL5A�JEC1��B�WA�ir����°�C��B����0��BI�$A﯇�	�.��y�E��(�B��L��
B�f���Q��B�� Bg��C��L       split_indices[$l#L       s      	               
      	   	                   
   
       
             
                                                   	                            
                                     
                                                                                                                                                                                                                              L       
split_type[$U#L       s                                                                                                      L       sum_hessian[$d#L       sE�8 E�p D�  E�� D.@ B�  DҠ E�P C� D  C  Bt  @�  C�  D�` C�� Eo� A�  C�  BP  C�  B�  B�  Bh  @@  ?�  @�  C8  C�  D�  A�  C�  A  B|  Ek� @�  A�  C�  B�  A�  B   C�  B�  BL  A�  B@  B  B0  A`  ?�  @   @�  ?�  B�  B�  C3  B�  D�  B@  A�  A   C"  C&  @�  @   A�  B   C�  ES� @�  ?�  @�  A   CF  C  BD  Bd  @@  A�  Ap  A�  B�  C�  A�  B`  @   BD  A   A�  @�  B0  A�  A   AP  A�  A  @�  @�  ?�  B�  A0  B�  @@  B�  B�  BT  B  D�� A�  A  B  @�  A   @�  @@  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       115L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       q?I60Au���"�BT����VV��X@Em�B���B��"����CU�������C`C��6��B�q�Bs|�C��C//�F�í�3�r�22pC�Bm�Z��]#7»(:Ë�SD���y� C	��¢�YC�bEA#*�B�#H�=�1C�d�䶑B��C�)��l���I������`K�p��l3�ǔ]C
�5B�3CV<�f�A�)��S���{��1	e�Õ��؍tC6�fB+�:B���9��R��C��+Ϝ���VC(,
�縉B��*��s��*�A�"�CI�ôRU�T�C�B�hR¼~A�DDc�A�A�C���C��dzë �%0YB'�m]#B��Q�u�9����A��RBa4%@�!��ׇ�B(H����Bmi@��:B����~H�A�/��4��iO��bA�������	IvBn������-A���ygL       
categories[$l#L       ?                      
                
                                   	   
                                            	   
                                                    	   
                   L       categories_nodes[$l#L                                   $   +   0   1   >L       categories_segments[$L#L                             	                                          +       ,       /       =       >L       categories_sizes[$L#L                                                                                                  L       default_left[$U#L       q                                                                                             L       idiL       left_children[$l#L       q               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W����   Y   [����   ]   _����   a   c   e   g   i����   k   m������������   o��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       qI�g�JD��I���J���JFYMI[��I�OlJ��J�HXJ�I[Jp{ I˯lI]�IDޘI"�J��J�s3J�t�J�� J��,JFUJ�/�J9H��I^��I�I�WI;�I"mG� G���J��fJ���K*��JG$&JSJDJ��J>��J�UOK\�GI���Ji@PI38    JU�!J-�k    FUxG�!�    I�HJ�Ie�tI>r�I �    H�*PIl��            F�                                                                                                                                                                                                        L       parents[$l#L       q���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   -   -   .   .   0   0   1   1   3   3   4   4   5   5   6   6   7   7   9   9   :   :   >   >L       right_children[$l#L       q               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X����   Z   \����   ^   `����   b   d   f   h   j����   l   n������������   p��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       q   @*=qB�aH>��>-V<#�
@o�P>�ZB�  @Å<���D��          =��m   B�     >��Bt  B�  >��
   B33D�� ?��?��?�bN   @�  B�  >	7L>���>���>�   @�  B�  A�  B�aH<�C�?�F   ��`K>bM�D�� �ǔ]      CV<@��HB��=?��FB  >\�1	e>49XB�  C6�fB+�:B�   �R��C��+Ϝ���VC(,
�縉B��*��s��*�A�"�CI�ôRU�T�C�B�hR¼~A�DDc�A�A�C���C��dzë �%0YB'�m]#B��Q�u�9����A��RBa4%@�!��ׇ�B(H����Bmi@��:B����~H�A�/��4��iO��bA�������	IvBn������-A���ygL       split_indices[$l#L       q                
         
                                      
                                              
                                    
                                 	                                                                                                                                                                                                                                 L       
split_type[$U#L       q                                                                                                    L       sum_hessian[$d#L       qE�8 E�� D�  EP EY� D�  B�  D�� DT@ C�� EHP Ap  D�  B�  A   D?@ D� D5  B�  CY  Bp  B  EF  @�  A  D<� D� B�  B  @@  @�  B�  D @ B�  C�  D3  A   B�  A�  C#  BX  B4  Ap  A�  @�  C  E<� @�  @   @�  @�  C�� C� C�  C  B�  @   A�  Ap  @   ?�  @   @@  B�  B8  A�  D@ B�  B$  B(  C�  C   D  @�  @�  @�  B�  @�  A�  C"  ?�  B  A�  @@  B(  @�  A  @�  A�  Ap  C  E*p C�� ?�  ?�  ?�  @@  C_  BP  C�  AP  C�� B�  BD  B�  B<  A�  @�  A�  A   @�  @   ?�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       113L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       u?օ�7W@�$��A��A�V�ϼA�&¡��B��W� fA_��i��*jZBȅ��5v�B����U�E���Bj�vC���{2B��X���BŠu�CZ�*��È�¡�5C�JBC*{�q5�A��C�/������~8����R�
C�+PAHV�C�ACz>]������O���>CCl@�B}��9�C�)oAʧ��k�+�k7�<��B�2��AҴ�&��ÿzkAë+A�K�D?t�¯ �A%L��^�nB��DC!����g�)4�B���.��M��A�����t�����H���aCW�+A���#�C�;A+��BT���K�A�N�.ܛ���*BT�B�Z�Ad�0�T$UA��U7���yAmA�Cڸ�@��(BA��A�w��k��ξ�¥"�©��BqR�BÒ?�.zB6��)Ç77�4*��5j�AA՚B��F���iB�n�UYoB��wC�e�L       
categories[$l#L       %                               	   
                   
                       	                                
          L       categories_nodes[$l#L       	                  "   '   ,   3L       categories_segments[$L#L       	                                                                $L       categories_sizes[$L#L       	                                                               L       default_left[$U#L       u                                                                                                     L       idiL       left_children[$l#L       u               	                                    !   #   %   '   )   +   -   /   1   3����   5   7   9   ;����   =   ?   A   C   E   G   I   K   M   O����   Q   S   U   W   Y   [   ]   _   a   c   e   g   i   k   m   o   q   s��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       uI�'�I�!dI�s�IN��IӟAI۾oI�#�I�#�I^�DI��I%�JɒJ�VI���Iؼ4H�I��IL�I�E~I��Ib�H�a�H���Jv�TJ��I�-
    I�k�Iǉ,I4�,J ��    H�M�IXF]Ie�H|��IS�I(d�I��I�g�I�IY�>    Hѫ�H��H��H�b�J2u1J��,K��J/�J*��I�#�I��I��I:	TIh�I{�H�I,IF��IO!(                                                                                                                                                                                                                                L       parents[$l#L       u���                                                           	   	   
   
                                                                                                                             !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <L       right_children[$l#L       u               
                                     "   $   &   (   *   ,   .   0   2   4����   6   8   :   <����   >   @   B   D   F   H   J   L   N   P����   R   T   V   X   Z   \   ^   `   b   d   f   h   j   l   n   p   r   t��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       uB     A&�\>+   ?(�9>���?p��   >�z�>���>�9XC  ?�ȴ   =q��@�  @i��D�� =o@j��D�  A��H@�  >�Q�   CZ�*>s�FB�
=?'+Bt  BC*{>V@߮   @_\)D�@ @@  >T��   @�  @�33Cz>]=�
=   ?��R>�=qA�  B�33B�  B|     @@  >Õ�>���=� �B�  A�  D�  >u@@  ¯ �A%L��^�nB��DC!����g�)4�B���.��M��A�����t�����H���aCW�+A���#�C�;A+��BT���K�A�N�.ܛ���*BT�B�Z�Ad�0�T$UA��U7���yAmA�Cڸ�@��(BA��A�w��k��ξ�¥"�©��BqR�BÒ?�.zB6��)Ç77�4*��5j�AA՚B��F���iB�n�UYoB��wC�e�L       split_indices[$l#L       u                                	                                                        	      
                                                                                                                                                                                                                                                                                                                                L       
split_type[$U#L       u                                                                                                            L       sum_hessian[$d#L       uE�8 Dt@ E�� D$� C�� E�� C  B�  D	� B�  CX  E�� C�� B�  B  A�  B�  C�� C)  B�  A�  C&  BH  E!� E; C�  @@  Bh  B`  A�  Ap  @@  A�  B�  A   C�� B�  B�  B�  A   B�  A�  @@  B�  B�  A�  A�  E  C�� Bt  E7@ Ci  C  B   A�  B@  A   @�  A�  A  @�  A�  @@  B�  @�  A  ?�  C  A@  BH  B�  A�  B(  B  B�  @@  @�  Bl  A�  A   A  A  B�  A`  B|  A�  @�  A0  A�  D9  D�� C�  B|  B@  AP  E. C  B�  B�  B�  BD  A�  @�  A0  Ap  @�  B,  @�  @@  @@  @   @�  A@  @@  @�  @@  @@  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       117L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       Y?�J�u�CM�@����2��Cێ!B��!@/��C1y���Akx�6C���Ï!�@r��D�VB���Co��_IcC�>����%B����<�C+P�DD,G�Bל�A�n4� E�C��C���C��C(._�p����>�D1��@�#�Òw�C������\P�Ì�uC���خ�C�o�B[�­��U�LB�:��A�{�$N��;�@<>B��i��@��{�D$�C!?QBI�A#�Cl�]V��C  ��6�N/�C�C£m�B���C�+��[���sZ5C�;�B����V�C��>��4�*�jB���A.u�§Y�C��i_mBI� �Pu�L       
categories[$l#L                                       	   
                                  
             L       categories_nodes[$l#L                   '   +L       categories_segments[$L#L                                           L       categories_sizes[$L#L                                          L       default_left[$U#L       Y                                                                              L       idiL       left_children[$l#L       Y               	����                                    !   #   %   '   )   +   -   /   1   3   5   7   9����   ;   =   ?   A   C   E   G   I   K   M   O   Q   S����   U   W������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       YI�xJI���J]ZJ
QJ#�
    IՏ\I�4J�JJ�J��J	��I�z�IЁ�Iө�JS�(I�:I��JT^J���J�&I�IAo�I��^H�@H�#�Ic��J\�I�3�I�Њ    I���I���I�g>I�\8J=hJg�\I��JE�DJ4�JH��Ha� InT�G�    IF@J��                                                                                                                                                                        L       parents[$l#L       Y���                                                     	   	   
   
                                                                                                                                   !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   -   -   .   .L       right_children[$l#L       Y               
����                                     "   $   &   (   *   ,   .   0   2   4   6   8   :����   <   >   @   B   D   F   H   J   L   N   P   R   T����   V   X������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       YA@  @�  =�hsC  >P�`Cێ!>���<49X=��
Bh  =�PB�     >L��   @�  ?°!=�wA�  B7��B�     >�7L>��B�  Bf  >>v�B�  >o��>���C��?M��D�@ B;��?z�<�`B?�(�@)��D�@    D�� B_�D�`    Ì�uD�� B�  C�o�B[�­��U�LB�:��A�{�$N��;�@<>B��i��@��{�D$�C!?QBI�A#�Cl�]V��C  ��6�N/�C�C£m�B���C�+��[���sZ5C�;�B����V�C��>��4�*�jB���A.u�§Y�C��i_mBI� �Pu�L       split_indices[$l#L       Y         
                                  	                                	               	   	       
                                                                                                                                                                                                                      L       
split_type[$U#L       Y                                                                                    L       sum_hessian[$d#L       YE�8 E�� B�  E� DM� ?�  B�  E�� B�  C�  C�  B0  B  A�  E� A`  Bp  C�  B�  A�  C�  B  @�  A�  @�  A`  @�  E` Ec� A  @�  B   A�  A�  Ci  B�  BX  A  A�  C�  A�  @�  A�  @�  @   A�  A`  @@  ?�  A  @�  @�  @@  E� A   D�@ E� @�  @�  A�  @�  A  A�  A�  @�  CD  B  @�  B�  A�  A�  @�  @   A`  @@  C�  @   @�  A�  @�  ?�  A�  A   ?�  @�  AP  @@  A   @�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       89L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       Q?�#�_]�?���è�����sBW���E��5�>�����W�B7��B�	V��$�B������¬�)���1�V���U�@��j��S)�EvXC|��}>Cé�B�5�d]>=~���]����?~�4�&�4B#�B�j�CLB@D,QX����CӉ���P��AG.C��Ç�Õ�MÆK��_^~B� 
���c��A>z��Z,��KAU�FZB��%�8��@�{(¯��B�Fv���CΤB���$�>��m���	eC�����x�C2ý0��;TsB>}���C��B��Ȧ��t�@�*�� U�C6�AO���&��1��B��L       
categories[$l#L                         L       categories_nodes[$l#L                      L       categories_segments[$L#L                                           L       categories_sizes[$L#L                                          L       default_left[$U#L       Q                                                                         L       idiL       left_children[$l#L       Q               	               ����               ������������   ����   !   #   %   '   )   +   -   /   1   3��������   5   7   9   ;   =   ?   A   C   E����   G����   I   K   M   O��������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       QI��Ie�I��
H�H�H2 AJW�*I��JHC�DHW�PG �    J�	sJ*��JRkJ
�G=Fv            D���    JE?JrU�J7gJZ��J��H��J�J�oF)��E#��        I���IAr�JS<Ju��J<:K5��J5uJ>2�I� �    F8|@    I�O�K+�)I���Jov                                                                                                                                L       parents[$l#L       Q���                                                           	   	                                                                                                   !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   +   +   -   -   .   .   /   /   0   0L       right_children[$l#L       Q               
               ����               ������������    ����   "   $   &   (   *   ,   .   0   2   4��������   6   8   :   <   >   @   B   D   F����   H����   J   L   N   P��������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       Q<�t�?4��   @@  D�  >��uD�  >�;d@u@�  B7��BX  Bճ3@�     @   ���1�V���U�@   �S)BH  >Ƨ�B�  >���   @@  B�  @@  B     ?~�4�&�4D�` @   B�  >��HB�  ?+�>r�!>�I�?1hsÇ�B!  ÆK�D�` B�33>���?�ĜA>z��Z,��KAU�FZB��%�8��@�{(¯��B�Fv���CΤB���$�>��m���	eC�����x�C2ý0��;TsB>}���C��B��Ȧ��t�@�*�� U�C6�AO���&��1��B��L       split_indices[$l#L       Q                  	      	                                                                                                           	                          
                                                                                                                                L       
split_type[$U#L       Q                                                                            L       sum_hessian[$d#L       QE�8 A�  E�x Ap  A  D�� E�  A   @�  @�  @@  C� D� C  E�� A   @   @@  @   @@  @@  C�  CA  D	@ A�  C	  @�  E�� D� @�  @�  ?�  @   C\  BP  C/  A�  D� Ap  Ap  A   C  ?�  @�  @   E�� C  C�� C�  @   @   @@  ?�  B<  C-  A   B(  B�  BL  @�  AP  D  A�  A   @�  A  @�  @�  @�  C  @�  ?�  @@  E  E"� B�  B  Ce  B�  C�  A   L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       81L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       k>��A����e A�,C -��N{�?��¦��A�F���9�C%U3�e�%C������@�B��^����3�B�Q���Δìb��:�SB��Dr7��B1,I�擷D - �B�����A�c��^�N]_��?�B�����N�J�KB���ü	��58_B(� ��ő��yCs�����D�ZO��o��k�C�q*�1y%B/vgCYs�A��C6c��eP�C�|�wO�BR�,�;`�@��¾�yB�J����YB�B@`�B�['��?�ã,2A�;fB�i��~��Æ��C�mT���Bb����C ��·�\C���Br�C!�ZCޘA� ���������BG�@C��x�IB�DBӲE�B�G?�U= ��C)BXg�A%b�1[Bk&�@�C��NA9u1�';$Bh}��ix�� �L       
categories[$l#L                                                 	   
                                              	   
         L       categories_nodes[$l#L                          .   7L       categories_segments[$L#L                                                         L       categories_sizes[$L#L                                          
              L       default_left[$U#L       k                                                                                               L       idiL       left_children[$l#L       k               	                                    !   #   %����   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C����   E   G   I   K����   M   O����   Q   S   U   W   Y����������������   [   ]   _   a   c   e   g   i����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       kI�+�J"`�I�2�J�J��\I隦JF�J'�oJ/�%I��vJ�KI��I�6�I^U�I�ôJ`��I�paJ�pJ�x    I"�J��pJFE8J�1J/1�He-�H���I~��IRl�JI�J��IzI�LI�x�J5N�    I���I�l:I��H�|�    Jͧ�J�F    HTz�I��JU*J9�nI�ɒ                H���Ix�G� I�^J�gLI��JYi[J3�b                                                                                                                                                                                        L       parents[$l#L       k���                                                           	   	   
   
                                                                                                                                   !   !   "   "   $   $   %   %   &   &   '   '   )   )   *   *   ,   ,   -   -   .   .   /   /   0   0   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <L       right_children[$l#L       k               
                                     "   $   &����   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D����   F   H   J   L����   N   P����   R   T   V   X   Z����������������   \   ^   `   b   d   f   h   j����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       k   B�     =��?&ffC     >�9XD�  =���B�  ?��   ?�^5@��B@�@�  <49X=��ìb�@�  >ȴ9@   BM�>��D�  ?f$�>o��=���   @�  =�+@���@@  B�  �J�KA (�=�+=��w>\��ő=��m>�I�����@@  >:^5   @�  ?bJB/vgCYs�A��@�  >�P   >�7L@�  @�  A�  A�  B�J����YB�B@`�B�['��?�ã,2A�;fB�i��~��Æ��C�mT���Bb����C ��·�\C���Br�C!�ZCޘA� ���������BG�@C��x�IB�DBӲE�B�G?�U= ��C)BXg�A%b�1[Bk&�@�C��NA9u1�';$Bh}��ix�� �L       split_indices[$l#L       k                        
      
      	                     	          
         
                      	                   	   	             
                                                 	                                                                                                                                                                                                    L       
split_type[$U#L       k                                                                                                    L       sum_hessian[$d#L       kE�8 D�` E�` D�  CR  DW  E�� C�  D�  AP  CE  DT  A@  C  E~  B�  C&  DI� D8� @   A0  C=  A   D4� B�  @�  @�  B�  B�  EJ� DN� BT  B  B�  B�  @@  DI  A�  D4@ @�  @�  Bx  B�  @   @�  C�  C�� A`  B�  @�  @   @�  ?�  @�  B�  @@  B|  D�� D�` C�  C�  @�  B8  B  @@  B�  A�  B�  @   D:� Bd  A`  @@  ?�  D4  @�  @   A�  B8  @�  B�  @   @�  B�  C�� B�  C  A0  @@  B|  B@  @�  @   A   Bp  ?�  @   A�  B  C�  D�  D�� D� C�� B�  C�  B  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       107L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       s>�Z��?��@Z:�ԛ�B`)*Cw��=suB�����=����C�C�D	�VB�^R�H@�B�#�s�C�{���C�3�@�N_���D�gB�B(B��Db�C��B�����E>���D4��Bk
(B�1Âp�D),C\§� Þ(nB�._Cb�QB���K?�K�����tCQ��D��]Ce:�ð�aCF_	�$�� gD�9uDMKA��@C!��ۗb���ì#�B����~%D�_�Bc�A)��D�B����fO!��:�@xC���B�64B=<`²u���e[���ݎ�{)�Bc����ABj�E��BC�n#�C(�C�ٶB���AX�qC#���RXC�UڴBU��䅿C�j�B�&tCQ= Bp��BQ>�����B�����:A����:B߱~�֨�A
9�Ol�C\�A�q��]B4��D"SC#BM�W��Ḃ�AH���<c�Be�RC�k�L       
categories[$l#L       2                            	   
                                                                 	   
                         	         
                        L       categories_nodes[$l#L                                !   $   '   (   ,   -   3   4   8L       categories_segments[$L#L                                                                       "       #       (       -       .       /       0       1L       categories_sizes[$L#L                                                                                                                       L       default_left[$U#L       s                                                                                                  L       idiL       left_children[$l#L       s               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I��������   K   M��������   O   Q   S   U����   W����   Y   [   ]   _   a   c   e   g   i   k   m   o   q����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       sI��JRJ�$J��JBrJ���J��I��vJ�I�NhJ��J��ZIel�J�J���IL>JcJ##�G���I��HG��Jq�I�r�JaWJtI%�Il4JH^�J��KҒJq�XIqH��nH��(H�6BI���J1
        I��3I��\        Ij�*H���I�p�H�"    I,o�    IZ� HG�A)IM��I)LJE��J��aJ���I�`&I�J�J6��J
zv                                                                                                                                                                                                                L       parents[$l#L       s���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   $   $   '   '   (   (   +   +   ,   ,   -   -   .   .   0   0   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <   =   =   >   >L       right_children[$l#L       s               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J��������   L   N��������   P   R   T   V����   X����   Z   \   ^   `   b   d   f   h   j   l   n   p   r����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       s?&ff>^5??:�H>%@@     B�  B4(�   ?Q&�B�  D�` D�  <ě�=�jB�\         B@�D�@ >�b>8Q�@@  B33>��y   B�aH=0 �>(��B�  =�^5      >�  @�     B�._Cb�Q      �K�����t=�1      @�  CF_	Bt  �� gB�ff      >V>)��=���   =��A@  @�  <�h@�  >��B����fO!��:�@xC���B�64B=<`²u���e[���ݎ�{)�Bc����ABj�E��BC�n#�C(�C�ٶB���AX�qC#���RXC�UڴBU��䅿C�j�B�&tCQ= Bp��BQ>�����B�����:A����:B߱~�֨�A
9�Ol�C\�A�q��]B4��D"SC#BM�W��Ḃ�AH���<c�Be�RC�k�L       split_indices[$l#L       s                                              
                                  
            	                                                                                   
      
      	                                                                                                                                                                                                                               L       
split_type[$U#L       s                                                                                                   L       sum_hessian[$d#L       sE�8 C�  E�� C�  C  B�  E� B  Cm  B�  B   A�  Bl  Eǘ C/  A�  A�  Ci  @�  B�  @�  AP  A�  A`  A�  A   BL  CI  E�P A`  C!  A0  A   A   A   C"  B�  @@  ?�  B�  A�  @@  ?�  A   @�  A�  @�  @�  A   @   A`  @�  @@  A�  A�  C  B4  C�  E�� @�  A  C  AP  @�  @�  @�  @@  @�  @�  @�  @�  B�  B   BP  A�  B,  B,  A   A�  @@  @�  @�  ?�  A`  @�  @�  ?�  @�  @�  A@  @   @@  @   ?�  @   A�  A   A0  AP  A�  C  A�  A�  A@  C�  E�� B|  @@  @   @   @�  C  @�  A   @�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       115L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       u?@�N�A"_i���5BѸ�)�NAG�ع.�e�wC�CC¨_oB 9�ƽ���
�BD���'�C����pd�4~|C<n{Dp,����{D3JC���Jŗ²"/�(��)�?���A���C���cY��s�A��&D`4�A�'M��!��O�C��U�LxeC�gD�q��q� ��I��[4�BMo�C������fC��Y�c@ �E�ÀX�C&�)Aj��\�n@���P�}��r�C��A7��C(Y5C��D�EW�6r�BV�@��`�J�`A��H��D YRB�fG�;AǶ|�xs(��Z��4B�@6CM��*@���e��B���f�TC�'�¤n�@�~g��ȷ�8l�B���A�nJ���z��� B�p�A��6�P�*�'aE�ݫ�`��B��m�3��ÎN[A����C��:MA�F�<��_�%��Ay��C$]@��C�@��Co,B��K7���i�D[%L       
categories[$l#L                                                     L       categories_nodes[$l#L                 !   (   *   1   5   6L       categories_segments[$L#L                                           	       
              L       categories_sizes[$L#L                                                               L       default_left[$U#L       u                                                                                                       L       idiL       left_children[$l#L       u               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W������������   Y   [   ]����   _����   a   c   e   g   i   k   m   o   q   s������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       uI^�J��I��
I���J�<�JhKIѰ>JE�J��AJ���J$|�I8�5I�*@I���J�|0J-pJǜI�g�Jw��J!�eJ��bI���ID;tH�@�H�u�I�ʘI��hI��I�T�J@��K*��I;�I��wH춟J��lI���I�J9dI�!`I׹[J"t�Jb��G�]JI���            G��8H\�`G��x    G�I8    H��0H�j�IaE9JI-I�I�I���JEP2J� J::�J���                                                                                                                                                                                                                        L       parents[$l#L       u���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   /   /   0   0   1   1   3   3   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <   =   =   >   >L       right_children[$l#L       u               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X������������   Z   \   ^����   `����   b   d   f   h   j   l   n   p   r   t������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       u>fffB�  <�`B>-VB�  BV  A�  >+Bf  >�bN?��\>A�7B  >�ƨ>޸R<���B|  >�ȴ?�?}   D�� ?@A�B�ff>?|�AP  <���<49XBb  C  B�Ǯ?z�?49X      @   >�K�>�l�@Nff?�\)?}p�   >C��   >�V�[4�BMo�C���D�  B\)   �E�@�Q�C&�)      @`B>�=qC  @@  AP  >�$�>�B.  �6r�BV�@��`�J�`A��H��D YRB�fG�;AǶ|�xs(��Z��4B�@6CM��*@���e��B���f�TC�'�¤n�@�~g��ȷ�8l�B���A�nJ���z��� B�p�A��6�P�*�'aE�ݫ�`��B��m�3��ÎN[A����C��:MA�F�<��_�%��Ay��C$]@��C�@��Co,B��K7���i�D[%L       split_indices[$l#L       u                                          
               
                                    	   	                
      
          	       	                                                             	                                                                                                                                                                                                                           L       
split_type[$U#L       u                                                                                                             L       sum_hessian[$d#L       uE�8 E8� E�� E/` C  BL  E~� D�� D\  B�  B�  A�  A�  E  D�  D�� B   D  C�  B�  A  B�  @@  A�  A   A@  A@  CD  E� D�  B�  A   D�� A�  A0  C� B�  C|  A@  AP  BT  @�  @   B�  @   @   ?�  A  A   @�  @@  A   @   @@  A  B�  B�  E� A�  D�� C  B�  @�  @�  ?�  D�� D6  A�  @�  @�  @�  C�  CU  B  B�  Cq  A0  @�  @�  A   @@  B0  A  @�  ?�  ?�  ?�  B�  @�  @@  @�  @   A   @�  ?�  @�  @�  @   ?�  ?�  A   B�  B  B4  A�  EP @�  A  A  D�  AP  B�  B8  B  B  @   @�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       117L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       k?��AЛ��u���(��B�Q��G �S�YhTC�PB�窿�֮��49B<k��8�rI�BnÞr)AХ�C���BY��Ɓ@������Cf��I�A2�/ò�������R�B�ƌ��e�я��]�ZBByj�I�C�)�C/8� ���nt���d�pљA��d�=�����BF3C����$�.�ɑD. �A����O������,Bʾ��}�@�]�B�z�@�v���A�(�B_ ��	�m��(�KF&B�0�A$�A�|X�HW�B�3�C��B��CEu@IJ����A�'�RxB�A �+,�A��B�0K2���A��¤��B�V������2(>@$C5�hB��9V!�#��Æ�����?�_BaA�C��Bsn���}��#�܅#B���U����s���C��D���c�L       
categories[$l#L       1                                                          	   
                                  	   
                                      	   
               L       categories_nodes[$l#L       
                      "   *   2   6L       categories_segments[$L#L       
                                           	              "       #       0L       categories_sizes[$L#L       
                                                                      L       default_left[$U#L       k                                                                                                L       idiL       left_children[$l#L       k               	         ����                           !   #   %   '   )   +   -   /   1   3   5   7����   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a��������   c   e   g   i��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       kIB��I��HIh�RJ5mJI���I�*�I��V    J��&J�(Iʃ�J�D-I�j�I��0H6�rI�pIĀ�J���J	��I��OI��`I��LJ)� JTkI���G��PH��H��    H�s�I ��IrhI�C�I��J�sJx�J-GJ-0I��(J,�eJ��Jhl\J5HNI�&�J"�bJ�|�IudI湎H��I�K�        H"�&GܺH�a�Ir�                                                                                                                                                                                                        L       parents[$l#L       k���                                                     	   	   
   
                                                                                                                                   !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   5   5   6   6   7   7   8   8L       right_children[$l#L       k               
         ����                            "   $   &   (   *   ,   .   0   2   4   6   8����   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b��������   d   f   h   j��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       k   <���?�I�?,��>�ƨ@��H      C�PB�  A�  @�  D�� @�  BR  >�  =���=��
?p��>uB�  D�� =��B_�D��    @��A (�   R�   >9X=�+@�     >P�`>z�HB�ǮBճ3>I�@,��>�7L   @�  @�  A@  ?�\)B4(�@@  B!     ��O����@�     ?�ȴ@�  B�z�@�v���A�(�B_ ��	�m��(�KF&B�0�A$�A�|X�HW�B�3�C��B��CEu@IJ����A�'�RxB�A �+,�A��B�0K2���A��¤��B�V������2(>@$C5�hB��9V!�#��Æ�����?�_BaA�C��Bsn���}��#�܅#B���U����s���C��D���c�L       split_indices[$l#L       k               	                                          	               	                                	          	   	                              
                                                                                                                                                                                                                                          L       
split_type[$U#L       k                                                                                                 L       sum_hessian[$d#L       kE�8 D�� E�� B8  Dz  E�X C&  B4  ?�  C�� D@ E�� C׀ B�  B4  A@  B  C�� B�  C�  C  E~  D�� CM  Cb  B�  A   A�  A�  ?�  A0  AP  A�  A�  C�  A�  B�  C  C�� C  A�  E  D�  Bh  D�@ B�  B�  A   CZ  @�  B�  @   @�  A�  @�  A@  A  @   A  @�  @�  ?�  A�  A�  @�  B�  C  A@  @�  B�  A   B�  @�  C�  Ap  B  B�  @�  A�  C� D�  D6� D}@ BL  @�  D�` B�  B�  @�  B�  A`  @@  @�  A�  CH  @@  ?�  A�  B�  A   A   @�  ?�  @�  @�  @@  @�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       107L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       m>������"@u���z�lB�=nB��m?ko*B�q"µ1�C�Y�Ac�C�#M�;���-�@Ԧ�� pC]��@��CG7�D�uCg%����[C�[�·3��^��BG~��ښ��l�n@XuK�YR�C�¬�@C*!j§!k§��ã<����eD$� �3jNC�,NC� �B�=qC����D% �B��@/8 çJÐ��C�eC*��9�
�
��CN�@����=AO�����PBrpA��p�4p�A���B��A��y�@/	>�����B�48Bx!��r�QBɭCp��B_D�qA��<�C �CCTA�c��<DLA2HC��eB�$0�eA^C&��Y�B#��A�{���+�$}0�+0�B����oi���B� "��s�t����R���aT��A/&��#�����B�bD��E��e��ª�L       
categories[$l#L       6                  
                                  	   
                                                	   
                                                     	   
      L       categories_nodes[$l#L                                   "   %   9L       categories_segments[$L#L                      	       
                                   %       (       )       *L       categories_sizes[$L#L              	                                                                      L       default_left[$U#L       m                                                                                               L       idiL       left_children[$l#L       m               	                                    !   #   %   '   )����   +   -   /   1   3   5����   7   9   ;   =   ?   A   C   E   G   I   K   M��������   O   Q   S   U   W   Y   [   ]   _   a   c����   e   g   i   k��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       mI9!�J'��I�WfI��JGK�J�=�I��/H�ۄI��bJ���I��J�8I�1�I�I��IL�H�oXJ"�$I�dKI,xbG�m�    I�ѷJ|��I!SI�
I���I��    I�HWI��uI� H��OH�*�G��I��AI�n,IF4�HZaHHz[PILl        H�R�Ii�J�2J��H��wHly�I��pH��IϬ�H�g�I�    I�'KI[��H��H���                                                                                                                                                                                                        L       parents[$l#L       m���                                                           	   	   
   
                                                                                                                             !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   7   7   8   8   9   9   :   :L       right_children[$l#L       m               
                                     "   $   &   (   *����   ,   .   0   2   4   6����   8   :   <   >   @   B   D   F   H   J   L   N��������   P   R   T   V   X   Z   \   ^   `   b   d����   f   h   j   l��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       m>���>��>�(�   =���=�Q�>��
>R�   @   D�     >N�?�y   =�j>��@j�HB�        Cg%�   @�  >�O�@�  @�  A�  �l�n?��@�  D��    D��    > Ĝ>��   @�  D�@ =q��C� �B�=q?r�!>gl�>9X=uD�@ =��w@@  >�5?@�  A�  B��{CN�?M�B�33   D�` PBrpA��p�4p�A���B��A��y�@/	>�����B�48Bx!��r�QBɭCp��B_D�qA��<�C �CCTA�c��<DLA2HC��eB�$0�eA^C&��Y�B#��A�{���+�$}0�+0�B����oi���B� "��s�t����R���aT��A/&��#�����B�bD��E��e��ª�L       split_indices[$l#L       m                                         	            	                                                                                       
      
         
                      	                                                                                                                                                                                                                  L       
split_type[$U#L       m                                                                                                  L       sum_hessian[$d#L       mE�8 D1@ E� D  C  CA  E� B�  C�  A�  B�  B�  B�  BX  E�X BX  B8  C�  B�  A�  @�  @   B�  B\  A�  B   B�  BH  @�  E�� A�  A�  B  B$  @�  C�� BT  B�  @@  A   A�  @@  ?�  A  B�  B  A�  A�  @�  B  @�  BP  A�  BD  ?�  E�p B�  AP  A0  @@  A�  A   A�  A�  A�  @@  @   B�  C@  BD  @�  AP  B�  ?�  @   @�  @�  @�  AP  @�  @�  B  B�  A�  A�  A@  @�  A  A  ?�  @�  A�  A0  @�  @   A  B,  A  AP  B(  @�  E�� D�` B�  A`  @@  A   @@  A   L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       109L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       s>ƝA=m�
"DAӫ��jc�'Wa��*6��mB%1������-'�C��P�lm~B� w��kA�Gv�˓GB^����;C�F�����Z��I���qj�CU�ý�*¤�A�{�D�����ܩ���CL�a���C�n B8aB��5Al>�+��B�.^�Bg(@�l�"eR��ZA�1�¦v��»�B �g�����Bl�B����?�D#�� e��BGeDk��5���q�C������A����]P�CO�B¥�̗ ��>C�A�A}�g@�M�Aҫi�˛B-�J��qrA�{f�B�<#��4��gB�7����*�j��LBЉ���A�C��$a±�]�������!��A�Q���B/���A���!B�M��
B/3�C��`Av����CR��¬��Bs�?A�8'C�o�A�.E��%�&Csc�CE�¼~DA�g8�hǙL       
categories[$l#L                              
                           L       categories_nodes[$l#L                          #   (L       categories_segments[$L#L                             	       
                     L       categories_sizes[$L#L                                                        L       default_left[$U#L       s                                                                                                      L       idiL       left_children[$l#L       s               	                                    !   #   %   '   )   +   -   /����   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K����   M   O   Q   S   U   W   Y��������   [   ]   _   a   c   e   g   i   k   m   o   q������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       sI24�JrqI�>{J��I���I�g�I���J �YI���Ie(I_�+I��qIU��JI��I��I�b J2��I�s�I�\�H4I^ͬIaZZH���HB��    I2��H�@J�J[I|I�eI��
J#�5IƳRI�Z�J~��I���J���I�ZI�{�    E&
PI��KIz�IR?�I�܅H"�H�m        I'�GE�0H�HK��J��J1�XH�I_J5&I���J>s�I���I�C�                                                                                                                                                                                                                        L       parents[$l#L       s���                                                           	   	   
   
                                                                                                                                   !   !   "   "   #   #   $   $   %   %   &   &   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <L       right_children[$l#L       s               
                                     "   $   &   (   *   ,   .   0����   2   4   6   8   :   <   >   @   B   D   F   H   J   L����   N   P   R   T   V   X   Z��������   \   ^   `   b   d   f   h   j   l   n   p   r������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       s      =]/@�  D�` @�  =�j   @�  D�@ @T��@@  >A�7B�  =,1@Q�7B�  Bl  Ap        =��>և+@@  CU�>{�m=T��=T��>B�\=�P=<jBnffD�@ Bu�R@�     D�  D�� A�  B�.^   @   B�  D�� ?I�^?@  ?��mB �g�D�` @J=q>l�DAP  A�  A0  >���=��@�  @�  @��
=P�`A����]P�CO�B¥�̗ ��>C�A�A}�g@�M�Aҫi�˛B-�J��qrA�{f�B�<#��4��gB�7����*�j��LBЉ���A�C��$a±�]�������!��A�Q���B/���A���!B�M��
B/3�C��`Av����CR��¬��Bs�?A�8'C�o�A�.E��%�&Csc�CE�¼~DA�g8�hǙL       split_indices[$l#L       s          
            
                                              	                                                                           
   	                                                                                                                                                                                                                                                                    L       
split_type[$U#L       s                                                                                                            L       sum_hessian[$d#L       sE�8 EC0 Ew@ E� D1  B8  Et` C�  D�  CG  C�� @�  B   B�  Eo  Cv  Ch  D  C�  A@  C;  C�  A�  @�  @   A�  A�  B�  A`  B�  Ej� CI  B4  C[  AP  D�� C�� C�  BX  A  @@  B(  C  B�  CЀ Ap  A   @   @   A�  @@  @�  AP  @�  B�  @�  A   BX  Ap  A0  Ej  C  Bp  @�  B   C5  B  @   A0  DV� C�  A0  C�  B�  CJ  B@  @�  ?�  @   @�  B  C  A0  @@  B�  C6  Ck  @   AP  @�  @   @   Ap  @   ?�  @@  @�  A@  ?�  @   @@  Bt  @�  @@  @@  @@  @�  A�  A�  A`  ?�  A  @   C6  E^� L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       115L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       {>�.
A�����ٚB�@�@�:���{&C7��ziA��"��B�z,��A^���6�C�\�A���ݕDL3���DA���x��	?C�I�A�G��
r��M-i��B1B[���xMB�cZD�TB*�A9��C�i=A��bØ?�C]
C˕l���C^��B$�C����/m��*��@�6�Cل�B�g^�u�3Cn���߁C�)���W����B����d4�rT�B|ą@59��5B��pQ�C�����CY��CA�,�AJ`�C��@�XA�Rb�03Ü�_1����B�,�B�h��h��B��i��&�B!���]��A-�B�0eAZ��C����W'��tj���������B��C(XB���
�sB���AV� �9�mفB�9����7�AP�b¤��Ã�_��@��C j3�P�t�=�/��@�����'�A���B��ʿ����I��¼����$B�xCV"1A�7�L       
categories[$l#L       2                    
                         	   
                                  	   
                                                             	   
         L       categories_nodes[$l#L       
                               "L       categories_segments[$L#L       
                                                  "       #       $       %L       categories_sizes[$L#L       
                     	                                                 L       default_left[$U#L       {                                                                                                          L       idiL       left_children[$l#L       {               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K����   M   O   Q   S   U   W   Y   [   ]   _   a   c   e����   g   i   k   m   o   q   s   u   w   y������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       {I4weI��I���Jq��I��JM��I�3rJɉJ�1�I�Ij�2I�iJ-tyJ%�"Ig��Jep|I$�J-yQJ
�TI��I�|I��~I�I�BI��BI͢ J��J^�dJ-IG��JjC�Jb�I�.I.�JH���I)OcJ8�G��t    I���H���J?(nI�sIz4I���I��H
WH��I2��IA��IFI]I��    JJQEBJ��J�5I�QJC!Ip�7Ii&�I�oJ%5                                                                                                                                                                                                                                                L       parents[$l#L       {���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   $   $   %   %   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <   =   =   >   >L       right_children[$l#L       {               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L����   N   P   R   T   V   X   Z   \   ^   `   b   d   f����   h   j   l   n   p   r   t   v   x   z������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       {   >:^5>��A�     =�/      >49X=� �?#�
>F��BnffD�  @�     B�        D�� =   ?o�D�` >��H@�  >��`>�bN   >["�@~{>�\)B  ?�   D�� <���A�  C˕l=�%?M��D�` A�  B2  =�O�D�  ?�O�>VA0  D�@ >'�@�  C�)�B��{B�  >�v�>׍P=��w?�w@�  B�  @�  >�A���CY��CA�,�AJ`�C��@�XA�Rb�03Ü�_1����B�,�B�h��h��B��i��&�B!���]��A-�B�0eAZ��C����W'��tj���������B��C(XB���
�sB���AV� �9�mفB�9����7�AP�b¤��Ã�_��@��C j3�P�t�=�/��@�����'�A���B��ʿ����I��¼����$B�xCV"1A�7�L       split_indices[$l#L       {                                       	                            	            	      	         	      
                          	   
                  	   	                                                                                                                                                                                                                                                                                              L       
split_type[$U#L       {                                                                                                                 L       sum_hessian[$d#L       {E�8 D�` E�` C�� D�@ D  E�� C%  B�  D�� C�� B�  C�  E,� D�� Bp  B�  B�  @�  B�  D�@ C  B�  B   Bh  C�  C  D�� D�  D�� B�  B,  A�  B�  @�  BT  B@  @�  @@  B�  Ap  C	  D�  AP  C  B�  A�  A�  A�  B(  A�  C�� ?�  B�  B4  C}  DP  D@ D�` D� D�� B�  A�  @�  B  @   Ap  B�  A0  @@  @   B  Ap  @�  B0  ?�  @@  @�  B�  A@  @@  B4  B�  D�� A�  @�  @�  A   C  B�  A�  A�  ?�  A0  A  A�  @�  A�  A@  @�  A   C�  A�  B8  B$  A   B  CZ  B  A   DM� B�  CԀ C�� DQ� AP  C�� D�  A@  B|  @�  A@  A�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       123L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       {>��r@�v�����a�dAzNt�yH?@²ֿ�Ə­!����A���˂�C_dBO=�C���.mD��,Y�m��A���
_���
BM		��Ô�C�����C+)hA����hYgC�s�@<V���7D:(|�<� ��?A�����S���?�i�C�E�u]��RB�J��)(LB��C�}@���%W��&L��k�ICMZDK�$�ZC�ܗB�ɺC�~A���A��å	��F�JA.��D/�@bK��-±՞�1POA�3���~7����YAK�j�#�#�"2��/'MA/B�j��C IB	N�� �����B���,ùC	C�@휬��ՅA���@�~�BFA>�B���B+����m��k%AX3�B	���İ��ٷ��4µ��B���B��(C��������"��C�y�� �>B��u��B>)�C��p��hA~k�������l� �X�:N�w_�3i�BH!��p�!C3aB�tL       
categories[$l#L                                              	   
                           L       categories_nodes[$l#L          	      "   +   .   1   :   ;L       categories_segments[$L#L                                                                L       categories_sizes[$L#L                                                               L       default_left[$U#L       {                                                                                                           L       idiL       left_children[$l#L       {               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A����   C   E   G   I����   K   M   O   Q   S   U   W   Y   [   ]   _   a   c   e   g   i   k   m   o   q   s   u   w   y������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       {I<6wI���I�=�I�ZDI��FJ�[JY�K`82J��{I��J�>JG� JkBI��I�4�I�`�K��Jk,LI���I.�PI+�JE�JvJ.�jJ���I�IÌGJ:u>I���I^�dI9YzIϔ�I�    HL#BJ%�VJZ��G�*    H��H�TH�s�Iz�<J�[J��J$�JZe�J�WI�/4J+UVJ%*|I���I�}�I��J �eI�YdJ�]~I��Ic�%Iw�2I_o�Ha�mGnH                                                                                                                                                                                                                                                 L       parents[$l#L       {���                                                           	   	   
   
                                                                                                                                         "   "   #   #   $   $   %   %   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <   =   =   >   >L       right_children[$l#L       {               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B����   D   F   H   J����   L   N   P   R   T   V   X   Z   \   ^   `   b   d   f   h   j   l   n   p   r   t   v   x   z������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       {@�  >'�?CS�B�  B33>���D�` B�  ?�o   A@  B�  ?�!   A�  @�G�@@  >D��@�  @�<���@�  ?�7>aG�A   @�  @�  A   A@  >hs@I�?+�?St�D:(|   @�  > Ĝ>�+���>���@   >�=q=o   D�  >���   D�� ? Ĝ   @�Q�>���D�  B�  @�  ?�"�D�` @�\)      =�C�?C�B�=q@bK��-±՞�1POA�3���~7����YAK�j�#�#�"2��/'MA/B�j��C IB	N�� �����B���,ùC	C�@휬��ՅA���@�~�BFA>�B���B+����m��k%AX3�B	���İ��ٷ��4µ��B���B��(C��������"��C�y�� �>B��u��B>)�C��p��hA~k�������l� �X�:N�w_�3i�BH!��p�!C3aB�tL       split_indices[$l#L       {         
                  
                                                                                         	             
                      	         	            
                   	                                                                                                                                                                                                                                                   L       
split_type[$U#L       {                                                                                                                   L       sum_hessian[$d#L       {E�8 E�0 D�  D�� Ek  D� Dd� D�� C�  D�� E(� C�  B�  C�� C�  D�  @�  C�� @�  C�  D:� D|� D�  Cŀ B�  B`  B  B�  C C�  A   D�@ C  @@  @   B�  C?  @�  ?�  C�  B  AP  D7@ C�  D8@ D�  C�  Ce  C&  Bp  A0  B,  AP  A�  @�  B�  A�  C�� A�  A0  Cŀ @�  @�  D�@ B�  B$  B�  ?�  ?�  A�  B@  C5  A   @   @   C'  B�  @   B   @�  @�  Ap  D3� B  Cm  D
  C9  D�� C  C*  C  B�  C  C  A�  A�  B  @�  @�  @�  B  @�  @�  A�  @�  @   @�  A�  B\  A�  A   BD  C�  A�  @�  @�  @�  A�  C�  @@  @   @�  ?�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       123L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       s>���A!u���G�A�V4��)�������Xd�VϰBA8%B���ܰk�2��B��BYg;�0�U@����w�5B~d5�*0xD4yB6~��k�<A�m��D�\��BZ
E�5�f�B�#���~�ìt2�<��Bu��Be�&�@B��BA���� ����Bhg�C�eC��x�:�F)���C�@t���*���0��(^á�C:A���C=h�5QB>:�s:��	��C���B��+��#H�Fڣ��c�@ʸ�B�dw�kþ��©Z�A�\�B���@;�4�2Aې�B1m���YB��[�����r�A9DHC
�'�=��W�!CW7AJ��CGY�A��Q�6r��NCʛ��e��H��{UU@�����	�AFkA�KB����e�gAG=QB���"����g���+��&�B_~���������@����C#)AM^�BQ����@4�x�k�j,�L       
categories[$l#L                           
               	                                
                               L       categories_nodes[$l#L                             -   5   7   9   ;L       categories_segments[$L#L                                                                                     L       categories_sizes[$L#L                                          
                                          L       default_left[$U#L       s                                                                                                      L       idiL       left_children[$l#L       s               	                                    !   #   %   '   )   +   -   /   1   3   5   7����   9   ;   =   ?   A   C   E   G   I������������   K   M   O   Q   S   U   W   Y   [   ]   _   a   c   e   g   i   k   m   o   q������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       sI'7I��IhzI��EI���Iu��IEu�J��I��JP	I���I�(*I�0�H�hI#�HI˩8J��wI�Z�IHe(I�\�I���I��I�h^I|*�H��I�M�I1-H�I    I2w�I	<I���JT�J/wlILwFIܪ�I��-I8ċ            I��^IFG�I��I�- H��I�(!I��I���Hk6�H%PI�{�I��yH3�I%�HusG�\I4F�G���FԐPIl��                                                                                                                                                                                                                        L       parents[$l#L       s���                                                           	   	   
   
                                                                                                                                   !   !   "   "   #   #   $   $   %   %   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <L       right_children[$l#L       s               
                                     "   $   &   (   *   ,   .   0   2   4   6   8����   :   <   >   @   B   D   F   H   J������������   L   N   P   R   T   V   X   Z   \   ^   `   b   d   f   h   j   l   n   p   r������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       s   ?Ix�@u�>A�7=�x�?��?~5?B�ff   =y�#??}?�hs   @�  B\33>ȴ9B�Ǯ@�  @�        Bp  =oA��   ?�"�>2-?�uB�#�@� �@��=��-B|  @@  D�� >�V>�;d@@  ���Bhg�C�e@�  D�` <�C�?�ff   ?N�A\)@�  D�� A   B\  ?�M�   BR     B
ff   B2     @�  �Fڣ��c�@ʸ�B�dw�kþ��©Z�A�\�B���@;�4�2Aې�B1m���YB��[�����r�A9DHC
�'�=��W�!CW7AJ��CGY�A��Q�6r��NCʛ��e��H��{UU@�����	�AFkA�KB����e�gAG=QB���"����g���+��&�B_~���������@����C#)AM^�BQ����@4�x�k�j,�L       split_indices[$l#L       s      
      	      
   
          	      	             
                                
             
                                                	                        
                                                                                                                                                                                                                                                 L       
split_type[$U#L       s                                                                                                        L       sum_hessian[$d#L       sE�8 EC0 Ew@ D�  D�` Erp B�  D� D�  B�  D�  EU C�  A�  Bd  D@ B(  D�` C6  @�  B�  D@ D  ER� B  Cր B$  A�  @@  B$  A�  C�� C�  A0  A�  D)@ C�  C2  @�  @@  @   Bt  B`  C�  C  @�  D � EN  B�  A�  A�  B�  C�  @�  B  A`  @@  B  @   @   A`  B�  CZ  Co  A�  @�  @�  A  A�  D� Bx  C�  C  A�  C  B  A�  A�  B  @�  C�  B�  @�  @   @@  CZ  C�� EM� @�  B�  A   A  A  A�  ?�  Bt  BP  A�  C�  @@  @@  A�  A  A   @�  @   ?�  A�  A�  ?�  ?�  ?�  ?�  A   @�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       115L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       {>k���L�A(�������pB�[� ��@�vÓ��B�@�AcA�0�B��t��YA�=`��yB;Cc�����K�&BI�H�S΃�p���^?C��XA��xCԮ�BPx[�����\;�ò��A#��έ�CT":�IV C�{B�w�ç���G�A�[	9A�+`C�m��rX���Í�eC.6D�\�i��VBhHC�

A�]�²YD��A�i/Cͩ?FO�� C��;�����$���;�4�0�UCT�q��"!�ZB�N��٤A����Z0C+V�B�D�Btr<½m��L��C�S�S-�Ê��A���t0K����B�pq�_\��E#�]��?�g����&�l�����k��@_L���SV©�#B�ҔCl��/#�@Ӱ�B�s�*�#D)CQM#�r�E�bauB�B�G\C��uBWp�.]���ʙB���AE�'C/��A��<�v���A��p ��H���>\:´�eA}��B�!�­�aC:o���gL       
categories[$l#L       0                         
             	                                   	   
                                        	   
                        	      L       categories_nodes[$l#L       	                      "   +   .L       categories_segments[$L#L       	               	       
                                   )       +L       categories_sizes[$L#L       	       	                                                        L       default_left[$U#L       {                                                                                                            L       idiL       left_children[$l#L       {               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I����   K   M   O   Q   S   U����   W   Y   [   ]   _   a   c   e   g   i   k   m   o   q   s   u   w   y������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       {I��I�uJ3��J(P�I�}6Jy�I��I��J�!7I�T�I�s�I�A>J�-InI�I�GxI'�
IL�;I���I�0IӃ�IVI���I�t�I.�I�v�I�� Ja*�I�M�I��KI���IT�1I/�SH� H=�G|l�I|�rIz�,    Hh; J �3J���E�� H@�VI�T    I���I�_XI-�I+��I�|KZ�JY�JZ��JE�J�4�Ib�I.��HǞ�H�� I�H���I"J�I�$R                                                                                                                                                                                                                                                L       parents[$l#L       {���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   $   $   &   &   '   '   (   (   )   )   *   *   +   +   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <   =   =   >   >L       right_children[$l#L       {               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J����   L   N   P   R   T   V����   X   Z   \   ^   `   b   d   f   h   j   l   n   p   r   t   v   x   z������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       {@�  <���   B\33>;dZB�  B�  ?<(�@�  >���>D��<o@�  B�  A�        D�@    B�  >�?�>�33>6E�B�  >���   B�  Bj��?���D�  ?%�T   >�V   >��D�  �G�AD�� B�  >�P=+>z�   C.6D?9X   BH  A   B�  AQ�@�  ?�{>�j@5B�  Bt  >`A�@@  @�  @�  >���>ٙ���"!�ZB�N��٤A����Z0C+V�B�D�Btr<½m��L��C�S�S-�Ê��A���t0K����B�pq�_\��E#�]��?�g����&�l�����k��@_L���SV©�#B�ҔCl��/#�@Ӱ�B�s�*�#D)CQM#�r�E�bauB�B�G\C��uBWp�.]���ʙB���AE�'C/��A��<�v���A��p ��H���>\:´�eA}��B�!�­�aC:o���gL       split_indices[$l#L       {                         
                                                                                                                                                                         
                                                                                                                                                                                                                                                   L       
split_type[$U#L       {                                                                                                                  L       sum_hessian[$d#L       {E�8 Ew� EB� B�  Eo� E p D�� B�  BH  D� EI� D�` Ct  D~� B4  Bh  A�  B  A@  D� A�  B  EG� A�  Dߠ B8  CF  Dx� A�  A�  A�  BL  @�  A   A  A�  A�  ?�  A0  C� B�  A   A�  B   ?�  B  EE` @�  Ap  D�  C  B  A   A�  C.  Dv@ A  A�  @�  A`  A   A0  A   A�  A�  @�  @@  @�  @@  @@  @�  A�  @�  @�  AP  ?�  A   C� @   B�  B@  @   @�  Ap  A   A`  A�  A�  @�  D�� D�� @@  @�  A@  @@  D�� A�  C
  @@  A�  A   @@  @�  A�  @�  B�  B�  Dt@ A   @�  @�  @�  AP  ?�  @@  A   @�  @@  @�  @   A  @@  @�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       123L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       m>/*�A�׳�C'���	*B�f�A������hA�=��3�ΠSB���?�ʬC:�5��z���ÁY�A��3Bˋ�����BF�'�c�C.�@�)�A���pE<C�\F��3�ù����@3e������[�ir�B=j�u�g�>�C[q�����C3#B�=\:�3�zB���C�Oo�E�B�z@���Cp��A��ÿ5OBg6�Dz*���Ó�q��MÍ��C���=6?7g�C�U��p�A��e@�ɀ�F�����Arc6B�&3������ ���B����4C�����Co����B���A�C�Q���{��®�P�}B8�B�3��A���C�~B��e�ہW�j1��{����oB���B��zC�%AB*���b�P²�B��AA�sB�?`Bu|����B�"�O�CffB�mW�U�=�"�b>�<uB��L       
categories[$l#L       %                      	                                        	   
                                     
            L       categories_nodes[$l#L                           "   /L       categories_segments[$L#L                                           
              L       categories_sizes[$L#L                                                        L       default_left[$U#L       m                                                                                               L       idiL       left_children[$l#L       m               	                                    !   #   %����   '   )   +   -   /   1   3   5   7   9   ;����   =   ?   A   C   E   G������������   I   K   M   O   Q   S   U   W   Y   [   ]����   _����   a   c   e   g   i   k������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       mHΥ�I���I��I��J<�JI^aCI*goI���Ir��J �I�}�Jcw�I�(I2i�H��I)��I���It6�    H-�J�rJp@�I���I��mJ�GII�cJ
O�I�9JC�/J4�    E^�#I��HᠼH�=�I��I7�            I뙒J�TI���I�h�I�%iJ:r�H���I���JJ!J�ݦH>�    I��    I3=�Jq�I�� I��:J=C�JG�                                                                                                                                                                                                L       parents[$l#L       m���                                                           	   	   
   
                                                                                                                             !   !   "   "   #   #   $   $   %   %   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   5   5   7   7   8   8   9   9   :   :   ;   ;   <   <L       right_children[$l#L       m               
                                     "   $   &����   (   *   ,   .   0   2   4   6   8   :   <����   >   @   B   D   F   H������������   J   L   N   P   R   T   V   X   Z   \   ^����   `����   b   d   f   h   j   l������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       m   Bb  =�E�BH  =]/B�  =ě�<o>VD�  >��PB�33>�ƨ>o��BnffD�` @�mD�  @"�BF�'A`  >�$�?�bND��    >z�H   @@     @�  >�Z���[   D��    A  >�n�>��7C3#B�=\:�3�z>�o>5?}>�z�>��=�FB_�   =49XD�� @�  >:^5Ó�q?+Í��BDp�>z�<�C�@   ?St�B   @�ɀ�F�����Arc6B�&3������ ���B����4C�����Co����B���A�C�Q���{��®�P�}B8�B�3��A���C�~B��e�ہW�j1��{����oB���B��zC�%AB*���b�P²�B��AA�sB�?`Bu|����B�"�O�CffB�mW�U�=�"�b>�<uB��L       split_indices[$l#L       m         	            	      
      	                        	                                       	                                          	      
                             
                                                                                                                                                                                                                      L       
split_type[$U#L       m                                                                                                      L       sum_hessian[$d#L       mE�8 D�� E�� D'  C�  C� E�� C� C9  A@  C�  C�  B�  B�  E�� A   C� B   C  @   A   C'  CG  C�� A�  B�  A   A�  B\  Ev� D�� @�  @   C�  B�  A  A�  C  ?�  @   A   B�  B�  B�  C  C�  A�  A0  A�  B   A�  @�  @   AP  @�  A�  A�  Eu@ A�  DQ� D1� ?�  ?�  A�  C�� @�  B�  @�  @   Ap  A   B,  B�  B�  B   A�  B$  B  A�  A�  B�  B�  C�� A�  @�  @�  @�  @�  Ap  A@  A�  A�  @�  ?�  @�  A   @�  A�  @�  A  A�  B�  Eo� @�  Ap  C�  C�  D#� B\  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       109L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       C>%2�@#���U?(�C[y��w��R�C���>��B�-
D|�yC}�4��T�ë�¸^0C; Z�/��>�� ��oC�,C���@g���
C����'�C\&zA�� � �2�?�2C0(��+�QC���G� B�Ó9�Dj5B]��X�C��9A#[��� �ό�AFsA�W�ˬA@u�"C��B3f�¥��BTuVC^��§p�B�Y���!A�$}�ˌ1��V-B�u�C�JH�.	�B��g�0(�������CA;�L       
categories[$l#L                                      	   
                           	          L       categories_nodes[$l#L          
             !   #L       categories_segments[$L#L                                                  L       categories_sizes[$L#L                                                 L       default_left[$U#L       C                                                            L       idi L       left_children[$l#L       C               	                        ��������   ��������         !��������   #   %   '����   )����   +   -   /   1   3   5   7   9   ;   =   ?   A��������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       CH��AI�YCJKr:IfQ�J��JV�I��I|q(I{�I��I�gdI�0�I���        Gn8�        I<�I��.I�0b        H�q6JO��I�_    DpS�    I��XI� =J��I���I�>�IHPIG-�GˠIU��H�KuI�)^J��                                                                                                        L       parents[$l#L       C���                                                           	   	   
   
                                                                                         !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (L       right_children[$l#L       C               
                        ��������   ��������          "��������   $   &   (����   *����   ,   .   0   2   4   6   8   :   <   >   @   B��������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       CB�  B�  @�D� ?�=�jB0  >��mD�@ ?0��   ?:�H@   �ë�   C; Z�/��>�33=@�@�  C���@g>o��>+? �C\&z   � D�  ?:�H?�      BH��   Bb  =���<���>ؓu>	7LA#[��� �ό�AFsA�W�ˬA@u�"C��B3f�¥��BTuVC^��§p�B�Y���!A�$}�ˌ1��V-B�u�C�JH�.	�B��g�0(�������CA;�L       split_indices[$l#L       C                  
      
                                                           	                                           	         	                                                                                                        L       
split_type[$U#L       C                                                             L       sum_hessian[$d#L       CE�8 E� D� E�8 B�  D � @�  @�  E�  B�  @�  A�  C�  @   @   @@  @�  @   E�� BT  B   @�  ?�  A  A�  C�  @   @   ?�  A�  E�  A�  B  A�  A0  @�  @�  @�  A   C�  A�  ?�  ?�  Ap  Ap  C_  E� A�  @@  A   A�  A@  A  @�  @�  @   @@  @@  ?�  @   @�  @�  @�  Cր B  A   A   L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       67L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       G>}��>��r�b����B�+fõR^Bޫ@2ҥ��D�CR����R\��+���B
�g��0 ��жBc�v��å�A�$^C���B�a�\��BR����CPi@c^?���C�Ǭ����B�D�C_+"�����PD �=<.Ce0��G=7A�*���u��+v@��f�tB�Ӱ����BͶB��P�ibC���BY����vh�B@����.��HךB�b����-���/gA�ƺB�o�CAml����@�dSA���C�#�����{��¤�NA���L       
categories[$l#L                               	   
             L       categories_nodes[$l#L                !L       categories_segments[$L#L                             L       categories_sizes[$L#L                            L       default_left[$U#L       G                                                                 L       idi!L       left_children[$l#L       G               	                  ����������������                  !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E��������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       GH�
H�^�Hs��H�+#I��E��F�6I[��I�
�I�`�I��.                I�b�J�I�T0I���H�y�IL��ItX�I���I�S)I�Jx�]I�TI�8 I�>�I��PG���HRXH�tF�� H`H���I��I)�Hɹ                                                                                                                                 L       parents[$l#L       G���                                                           	   	   
   
                                                                                                                 !   !   "   "   #   #   $   $   %   %   &   &L       right_children[$l#L       G               
                  ����������������                   "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F��������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       GA��A@     A   >)��A���Bj��@�  B�  >o>�bN��+���B
�g��0 =e`B@�  B�  A   >�D�� ?"J>� �   ?M�=�1>�A�=��wA�  A   C  >B�\Ap     >L��>cS�A�  B\33=���A�*���u��+v@��f�tB�Ӱ����BͶB��P�ibC���BY����vh�B@����.��HךB�b����-���/gA�ƺB�o�CAml����@�dSA���C�#�����{��¤�NA���L       split_indices[$l#L       G                                                                                	         
            
         	                                                                                                                                            L       
split_type[$U#L       G                                                                    L       sum_hessian[$d#L       GE�8 E� @�  Eڐ B�  @�  @   E�� DW  B   B<  ?�  @@  ?�  ?�  E�H DK@ DR� A�  A�  A`  A�  A�  D5� E�� CA  D  DN� Ap  AP  @�  @�  A0  @@  A0  @�  A�  @�  Ap  C�  C�  EX� D�@ BD  C  C�  B�  A�  DI  @@  A@  A   @�  @�  ?�  @   @�  @@  A   @   ?�  @�  @�  @@  @�  AP  @�  @   @@  @�  A   L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       71L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       k>1Ƈ��}'@*]4�g(sB;Si�T>�@��Cd�$�C�WWA�¥�|��Ñ'DB��*@R��B��C鴬�J�G�s�!�Cp5��	�oD	E�a���x�C�x`�x(B|�?�IB�B'�dB���C}��UWCZ�(C��Í��©��B�M�D,��B�u�� Éa7CahB�����C!� �v6A�� ����C�Nê HCq�
B��p��s�5@�@sl�B~���)��B-�s� � Ak���*B�C�6*Bˮ\�����7���J�j�B��A�`BzB?���a� C���BD�5�Q����=BG A]���*�B9'�f����1��B���@�� ���4�M��B0v���$��pB���R�B�b�C���y&�Î��B�/�ﲭA���D	M�B&��&��qs¡�zA�I?�L       
categories[$l#L                                                            	            L       categories_nodes[$l#L       	      !   (   ,   -   .   0   4   6L       categories_segments[$L#L       	                      	                                          L       categories_sizes[$L#L       	                                                               L       default_left[$U#L       k                                                                                                L       idi"L       left_children[$l#L       k               	            ����                        !   #   %   '   )   +   -   /   1   3   5   7����   9   ;����   =   ?   A   C   E   G   I   K   M   O����   Q   S   U   W   Y   [   ]   _   a   c   e   g   i��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       kH��I�^OI'�\I��J<|�I�t�I7�II�I�U    I��I��I�Y�J�heI0�H��xI�f'I�LuJzI�!�I�6�I��$H�H��Ig,�J��'I��{J�I'�2    H>#G��    I�8pI��J��J@8I+��I�h1IӛH�9I?�'I.2    F�5�G8U�Gp�I�GX	-H���J�<VI�`�HZS�J�� I�ϩI���I��`                                                                                                                                                                                                        L       parents[$l#L       k���                                                           
   
                                                                                                                           !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8L       right_children[$l#L       k               
            ����                         "   $   &   (   *   ,   .   0   2   4   6   8����   :   <����   >   @   B   D   F   H   J   L   N   P����   R   T   V   X   Z   \   ^   `   b   d   f   h   j��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       k>��@e=]/D�  @j�HB�33>%�TB[��B�33C�WW>���B�  =�P>߾w=��   >["�B�  =��D�` =e`B=T��A   @�  B�  =���A@  ?ƨ=���B�B'A�  @�  C}�   @#�
>C�=�jB�  A0  >�\)   ? Ĝ>%Cah         @@     B\33>��B�     ?	�^   B�ff=�;dB~���)��B-�s� � Ak���*B�C�6*Bˮ\�����7���J�j�B��A�`BzB?���a� C���BD�5�Q����=BG A]���*�B9'�f����1��B���@�� ���4�M��B0v���$��pB���R�B�b�C���y&�Î��B�/�ﲭA���D	M�B&��&��qs¡�zA�I?�L       split_indices[$l#L       k   
                  
                                                                                           
   
         	       	                                                                                                                                                                                                                                                           L       
split_type[$U#L       k                                                                                                  L       sum_hessian[$d#L       kE�8 D� E� C�  C(  CU  E�` A�  Cƀ ?�  C'  C9  A�  B�  E�� A   @�  C�� B�  C  A�  C4  @�  AP  Ap  B\  A�  CB  E�� @   A   @�  @@  C�� A�  A�  B�  B�  Bl  @�  A�  C  A�  @@  @   A  @�  A@  @@  A�  B  A�  @�  C  B$  C�� E�h ?�  @�  @   @   B�  C8  A�  @   AP  @�  A�  B<  B�  @�  A0  B@  @   @@  A�  @@  C  A�  @�  A�  ?�  ?�  @�  @�  @   @   @   A   ?�  @   AP  @�  A�  @�  A�  @@  @@  ?�  C  ?�  A@  A�  C�� A�  B�  E�� L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       107L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       w>�2�A(���_�A����tA�3�z	YA���C��z�q�{�+���q��B,��A�߿�Ľ_B �.�WU¬D+VRCAγ��[������6��B ���	B�Ԏ�F��BL���c$¨�j���A��OC<��B}P��T3�A0��JC˵�C�P=D.�YB�BV��$�A�����5�]��A�W�!I�CÜ��ݤâ����C~
�BI�;Bk1�Lzw�7tB��÷[�@�l�@�����^C���i�[A�����(B�Cj9BgHh@�R|�9/���5�A���.��C�h@���A�6�Cw����B�&�D��B)�A��$�,�B]��Ob ���CC4ʝ�^�1Bo%���;B!\��3���BySB9���	z`B�VC9$g�/w\B �@�eB����*^�¥�B���e�C;��A�o�@�{M�	{6B"ug�A�����b��K1�B��!A��CAu�����ZL       
categories[$l#L                 
             	   
                           	   
          
                              L       categories_nodes[$l#L                                      #   'L       categories_segments[$L#L                                           
                                          L       categories_sizes[$L#L                                                                                    L       default_left[$U#L       w                                                                                                    L       idi#L       left_children[$l#L       w               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G����   I����   K   M   O   Q   S����   U����   W   Y   [   ]   _   a   c   e   g   i   k   m   o   q   s   u��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       wH�1-IF	IIt�I�i�I��hI�= I�!I�g;Jm�Ir��J-�I��@J-�J_J�tI��KI�AH I�IS-�I¹uIr9�I��I�Is�I�I�J0L I6�HJ��I�ŧJ"��IԺPI�[TI�A�I�;!I���E���    H�(    H�=�IBOI���I�h�HU    I/^    H�?�H��;I�BI/+zJ���JN��I��I8۹J!FJaN�I_g�I�*�I}�&JH��IŻ6I܈�                                                                                                                                                                                                                                L       parents[$l#L       w���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   %   %   '   '   (   (   )   )   *   *   +   +   -   -   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <   =   =   >   >L       right_children[$l#L       w               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H����   J����   L   N   P   R   T����   V����   X   Z   \   ^   `   b   d   f   h   j   l   n   p   r   t   v��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       w   ?>5?@�  ?<�      =Y�>߾wBH��=y�#?���      A  =Ƨ�>�t�         =�`B??}?��Bu�R?��>���>��D�  <���>��   D�` >H�9@�?�(�>7K�   �JB�33C�P=   @��
@�?}D�` D�� �]��Bt  �!I�>t�B�  B\33>�ƨB�  D�� ?s�F?pbN=�F=��>�(�>�;d@�  D�� ?�ĜD�  A�����(B�Cj9BgHh@�R|�9/���5�A���.��C�h@���A�6�Cw����B�&�D��B)�A��$�,�B]��Ob ���CC4ʝ�^�1Bo%���;B!\��3���BySB9���	z`B�VC9$g�/w\B �@�eB����*^�¥�B���e�C;��A�o�@�{M�	{6B"ug�A�����b��K1�B��!A��CAu�����ZL       split_indices[$l#L       w      
      
                   	   
                                                                            	                                                     
            	      	      	         
                                                                                                                                                                                                                                   L       
split_type[$U#L       w                                                                                                            L       sum_hessian[$d#L       wE�8 EC0 Ew@ D�@ D�  Dv  E9� D݀ A`  D�� B4  CQ  DA� D � E� D�@ D"� @�  @�  A�  D�� A`  A�  B�  B�  C�  C�� C�  Bl  D   D�  D�  B�  C]  Cր @�  @   @�  ?�  @�  A�  D8@ D� @�  A  A�  ?�  B   B�  B  B�  B�  C�  C(  CY  C"  C�  A�  B  CK  C�� B�  D�` D-  C�� B\  A   Bh  C#  B�  C�� @�  ?�  @�  ?�  ?�  @@  A@  A   D.� B  C�� Cf  @   @@  A�  ?�  @�  A�  Bp  Ap  A�  A0  A0  Bd  B�  A�  B�  Ci  C!  @�  CL  AP  A�  C  A@  C�  @�  A�  A�  A@  B�  B�  C�  A�  B�  @�  C0  D�` L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       119L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       {>�e2@�O��z���AE�^@����GP��Z��PE��s4A����w�QBX$C����)ޖ���^B�n�CG���W�M�Ao�wB���@�i��"��]�B����<©�B�G�_d"�����q2*��v�A3�1DL��M�C����l��w�@���[�+�8C\�Ϳ� �B����h��C�(����h�}F�kj��6��Ý�B&�!C��\�RJ�A���@�i�)�vC��~A�ؘ�I��>.i��79B��u�!BdB���C-���xB�=��K�"A��CCɜ�����AŐC,�M@�Y B��p�X����>�4#�t������ω����DC6K�A�qE@ÌS��F@�4�BL"�����A��UC���Z�A�x���hB?�G���v��)��}�*A�=���R@�ʈh� m�B�f=C�B9����h������B���£$�Aom�A�}���9y�C<�fB�'��5B%��x�0BN�S��L       
categories[$l#L                    
                            
L       categories_nodes[$l#L                    #   %   0   <L       categories_segments[$L#L                                                         	L       categories_sizes[$L#L                                                        L       default_left[$U#L       {                                                                                                                L       idi$L       left_children[$l#L       {               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c   e   g   i   k   m   o   q   s   u����   w   y����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       {H���I
�IPܞIRR�I�_�I\�I&�$I��)J���I.>I�\VH��"I8�I $I E�IɐFJ���J�*�J���IZŘI��J1�~J�TH��Hr�4INcJH��
H�3�I:XH��PIs�IxE�I��JvKPI���J5�XJE-�J �UId?�I0�I�^I LJ�I�]J�j�I��\H9�Fw1 F�afF�c�I��I0HR�H��H�-Hk}�H�D�H�4    Hp��Hoi�                                                                                                                                                                                                                                                    L       parents[$l#L       {���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   :   :   <   <   =   =L       right_children[$l#L       {               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d   f   h   j   l   n   p   r   t   v����   x   z����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       {   @�  D�� B�  B,  >�(�>�M�B�  >�7LA   @�  ?�ĜB\33   >���B�  @�  ?aG�>�1@�D�@    D�  >��T=ix�@+�B|  >?|�=�O�>���Bt  B�
=D�� @�  D��    D�     @�  >�v�>�B�\A�  A@  ?��F>333@�=��
   B8Q�@   B(  >�1'@�  @�  =��=�C�BV  ?��I�   >�\)B��u�!BdB���C-���xB�=��K�"A��CCɜ�����AŐC,�M@�Y B��p�X����>�4#�t������ω����DC6K�A�qE@ÌS��F@�4�BL"�����A��UC���Z�A�x���hB?�G���v��)��}�*A�=���R@�ʈh� m�B�f=C�B9����h������B���£$�Aom�A�}���9y�C<�fB�'��5B%��x�0BN�S��L       split_indices[$l#L       {                      	               
                                                      	                                                                      	                                                                                                                                                                                                                                                                                 L       
split_type[$U#L       {                                                                                                                    L       sum_hessian[$d#L       {E�8 E�p C�� El` E:� CA  B�  EUp C�� D�� D�` B�  B�  B`  B�  EG` Ca  Bl  C�  D6@ C�  DO� D�� B�  A@  B�  B   B  A�  B<  A�  E<� C)  CG  A�  A�  B$  A�  C�� D*� B<  A�  C�  C�  C�  A�  D�  Bt  @�  @�  A   Bt  A�  AP  A�  A�  A�  @@  Ap  @�  B,  A`  @@  E<  A0  @�  C%  B  C   A�  A   A   A   A�  Ap  @�  A�  Cb  Bl  B�  D� Ap  B   @�  A�  C|  B�  C)  C�� C*  C<  A   AP  C�� D3� @�  B`  ?�  @�  @@  ?�  ?�  @�  BH  A0  @�  A�  A   @@  AP  @�  @   A�  @@  A�  ?�  @   @   AP  @   B$  @@  A0  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       123L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       w>�����@���?X���A�4�F(BB#�o�X�C�B�����@8B�i�B=/��O����?i�I�=��C�B	k�D"eZ���C+�I��zBj�a�@	5SB�<C�=��������a�C2^�CG{Ô<fBr=���4DV��C
��C$ .��C��CVi�.�'�k�z����C�W�B���¿CB���?b�Cb�r�t��CF���mO0B�'u@�_�D{j�C"�E��CB��<�?��hC�XBu��C-`��ɧ��o�8^�B��v�>uyÐ3DB��fC���CP����CP���_A��J~>B���&�§�@'���cA���A����o��ի�CO���B���@���[A��B�y�B�B����
EB�W����EA:*K@�JoCˤ���sBx�
A�6�Cx�AS[����C�O#BT����%�B�aJ��FS�Cr?ZC�L       
categories[$l#L                                                                            	   
      L       categories_nodes[$l#L                !   "   *   0   9L       categories_segments[$L#L                                                         L       categories_sizes[$L#L                                                        L       default_left[$U#L       w                                                                                                              L       idi%L       left_children[$l#L       w               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9����   ;   =   ?   A   C   E   G   I   K   M   O����   Q   S   U   W   Y   [   ]   _   a   c   e   g   i   k   m   o   q   s   u����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       wH�l�I���I�^`I��7Jf�LI���I�v;I�ֹJ�gJ���J��Ij�BI�o�JZ�JZ�bI�X�I���I�u�J��4I�&�J��
JJ9�J3�I���I���IFa�I\�I���JcY    I2��I�:cJn��Ix�4I���I��#I��VJ=�JF{J\�I�FW    I5K!Jn�JF�JA�J'
I��I�)I��4J|�H]��I@lI�U�Ia4:J(O�I�I�x�I�0�H��H��'                                                                                                                                                                                                                                        L       parents[$l#L       w���                                                           	   	   
   
                                                                                                                                   !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <L       right_children[$l#L       w               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :����   <   >   @   B   D   F   H   J   L   N   P����   R   T   V   X   Z   \   ^   `   b   d   f   h   j   l   n   p   r   t   v����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       w?	x�B�  A�  B�  >�7LD�� ?2-B�aH@�  >��jA0  >'�>Q�?+?3t�?#o   >ɺ^=��>&�y=�^5   >;dZ>/�>�?}<�`B=�9X=��P=�C�����>P�`?`B=���      >x��B�  D�� Ap  B  D�  C��   ?�\>x��>�RB�  >N�   B�ffAp  A�  D�� B@  B�  B�  B      A�  =�\)?9X<�?��hC�XBu��C-`��ɧ��o�8^�B��v�>uyÐ3DB��fC���CP����CP���_A��J~>B���&�§�@'���cA���A����o��ի�CO���B���@���[A��B�y�B�B����
EB�W����EA:*K@�JoCˤ���sBx�
A�6�Cx�AS[����C�O#BT����%�B�aJ��FS�Cr?ZC�L       split_indices[$l#L       w   
                                                            	            	                      
            	                             
         	                                                                                                                                                                                                                                                                                 L       
split_type[$U#L       w                                                                                                                L       sum_hessian[$d#L       wE�8 E[@ E_0 E8@ D  E(0 D\  E3@ B�  C  C�  D@ E� DV� A�  E0� B,  B  B8  C  A@  C�  BP  C  C�  D� D�  DJ  BL  ?�  A�  E-� BD  A   B  A�  A@  AP  B  B|  B�  @�  A   C:  C.  A�  A�  B  B�  Ci  Ci  A  D@ A�  D�@ C�  D  @�  B8  A`  @�  E(� B�  ?�  B@  @�  @@  A�  A�  A`  A   A  @@  @�  @�  @�  A�  A�  B$  B  B  @�  @�  B  C  B�  B�  A�  @�  @�  A�  A0  A�  BT  B0  CS  A�  CS  A�  ?�  A   D  B�  Ap  @�  D�� A�  C�  @�  C�� C7  @@  @   A@  B  @@  A0  @   @�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       119L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       u?{?�^p�;,p���B5}]Bʯ�½u@�c��-$B�<F�ZECk���ԁ�ô�+�/\��G}?AźuA�����'h@���CJ�CJ?����C����}@B�k�×��V2?x���E�ä��C'5����SB^)�@�ׯB)'��@'�+��B��g�BW1�C�ݳ�{sCâĈg��x���@C�'gA�� �"V�C�{�4��b}���Ä�5�{JB����_CJ~�ö���EvB�kA�1(��`n�}�;@���B<�'��qh@˾�@���Bɔ�����Ð�1��7�C!��wF�r�Z3A��:��5Má�&�B)�B�ܱB���C�F���B��
¶kûؾ����b�A��{`A� �C/�An_� S4��� �o�gB��_A���0�W��A���	�ª#ç
���MB���A�����B�HK±���OI4���L       
categories[$l#L                                            
                              L       categories_nodes[$l#L                      (   -   /   1   3   8   9L       categories_segments[$L#L                                                                                     L       categories_sizes[$L#L                                   
                                                 L       default_left[$U#L       u                                                                                                        L       idi&L       left_children[$l#L       u               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W����   Y   [   ]   _   a   c   e��������   g   i   k   m����   o   q   s����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       uH��I��I��H�7�J,�lI��CIđJI�fqI���J�<J!k-Ir�^I�I݅2I-j_I��I�noJ1C�Ic`J���J@�XJ5�J
֬I|BxGp�@HKH��I���Hr?Iw��G�UXI��>I���J)��I�k�JDʺI�IbI��AI�F�J[I&s�J�Ji^ I.��    G�� H�<�G��CH�B D�i�E@� G�6�        G"i�I�wG�� H!;�    I��eI�W�G�p                                                                                                                                                                                                                            L       parents[$l#L       u���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   -   -   .   .   /   /   0   0   1   1   2   2   3   3   6   6   7   7   8   8   9   9   ;   ;   <   <   =   =L       right_children[$l#L       u               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X����   Z   \   ^   `   b   d   f��������   h   j   l   n����   p   r   t����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       u@�  B�=q>\)   >�VB(  >8Q�      >�~�D�� >:^5=D��B�  @?
=@   >�ffB�Ǯ@@  >޸RD�@ D�` >� �=@�@�  >L��B̊=>w��@�  ?ZD��    >�"�>�\)?�hB�  >��AP  B��{A�     >�7L>["�D�  Câ   @��   A�     B�     �4��b}�=ȴ9>��      �?WK�D�  @   �EvB�kA�1(��`n�}�;@���B<�'��qh@˾�@���Bɔ�����Ð�1��7�C!��wF�r�Z3A��:��5Má�&�B)�B�ܱB���C�F���B��
¶kûؾ����b�A��{`A� �C/�An_� S4��� �o�gB��_A���0�W��A���	�ª#ç
���MB���A�����B�HK±���OI4���L       split_indices[$l#L       u                              
                     
         
                  	      	                
      
                                                                  
                                                                                                                                                                                                                                                   L       
split_type[$U#L       u                                                                                                          L       sum_hessian[$d#L       uE�8 E�P C  E�� C�  B  B�  Ez� E"� C�� B  A�  Ap  A�  B�  D�� D�@ D+� D�  C%  B�  A   A�  A�  @�  A   @�  A   A   B�  @�  B\  D� D?� D�� D*  @�  D>  D�  C   @�  Bp  B(  A  ?�  @@  A�  @�  AP  @   @�  @�  @   ?�  @�  @�  @�  @�  @   B�  A�  @�  ?�  A�  B  C�  D�  D  CF  C3  D�  D!� B  @@  @@  D=  @�  D�� B�  A�  C  ?�  @�  A�  B  B   A   @�  @@  ?�  @   A   A`  @@  ?�  @@  A   ?�  ?�  @   @   @@  @@  @   @�  @@  @@  ?�  @@  @@  @@  B@  A�  AP  @@  ?�  @�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       117L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       e>o�RAq33�O�.A��6�5_�����@_ B��"���A�R�P8�C��A����?{���m9Cܰ�B�k��-�szA�6����1CH�п��d�8	Cqu��N%�)�B��.Ê|�k;[����C@.(D<��È�pC�H�B�9��vk��?�y(u�`�C�����~�����ȋC�An�I�
�i��?��Î�3���JC�9��=A�7T�c��BW� ¢���"��'����B��B���C����k��¾mA�_�C��B38@|�B%t������BՅ6®������B�)DB�AMFa�N��B����$��B�pGßЏC��c��@��>�;�A�c��G��TkB`͛�_���$C4��:B���C�<�B���/ �?ӯ�B��07�L       
categories[$l#L       '                                   	   
                               	   
                                         	   
       L       categories_nodes[$l#L       	               "   ,   .   /   7L       categories_segments[$L#L       	                                                                &L       categories_sizes[$L#L       	                                                               L       default_left[$U#L       e                                                                                        L       idi'L       left_children[$l#L       e               	                                    !   #   %   '   )   +   -   /   1   3   5   7������������   9   ;   =   ?   A   C   E����   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a��������   c������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       eH�� I��\J-�I���I��6IW�Jx�J(a�I�E*I1M�I�b�I�>�J0�7I �I�I�s�JL�I��I({I)f<H�ApIM�PIT��I(?�IMI�J*>I$n�H��            IZ>�I�{I���GJa(*I:� I��    Ii߂Ig�Fr�H}��I D�I�s�I��G�(I�3�ISFI+ͨI��JG26IH(�        F���                                                                                                                                                                                    L       parents[$l#L       e���                                                           	   	   
   
                                                                                                                       !   !   "   "   #   #   $   $   %   %   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   7   7L       right_children[$l#L       e               
                                     "   $   &   (   *   ,   .   0   2   4   6   8������������   :   <   >   @   B   D   F����   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b��������   d������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       e?���>F��B�  =�{>�?}B�  >�dZ?�z�>���?��R@�  Bd  ?�@@  > Ĝ?��      B�  >z�H>O�B�     >o��>�RD��    =�v�B��.Ê|�k;[?Y�B  >��\   >z�H>���@�  ��?>t�j>o��B(G�>�\)>ɺ^   ?+C�      B\  B�  @�  >>v�=� �A�7T�c��   ¢���"��'����B��B���C����k��¾mA�_�C��B38@|�B%t������BՅ6®������B�)DB�AMFa�N��B����$��B�pGßЏC��c��@��>�;�A�c��G��TkB`͛�_���$C4��:B���C�<�B���/ �?ӯ�B��07�L       split_indices[$l#L       e                                       
      	                                                                         
             	                                                                                                                                                                                                                                    L       
split_type[$U#L       e                                                                                            L       sum_hessian[$d#L       eE�8 D�  E�0 D�� C�� E�� A`  D)� C�  C	  C  E�� B  @�  @�  D&@ AP  C�� B�  B�  A�  B�  A�  E�  BD  B  @�  @�  @   @�  @   D  B  A  @�  B�  CY  B�  @@  BH  Bh  @�  A�  B�  @   A�  A  CM  E�� A�  A�  A�  AP  ?�  @@  @   @@  D@ B\  @�  A�  @�  @�  ?�  @@  B   A�  B�  B�  A�  B�  B8  @�  B  A�  @   @   A�  @�  A0  B�  ?�  ?�  A@  @�  @�  @@  BP  C  E� A�  A�  @�  A�  @@  A  AP  @   A0  ?�  ?�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       101L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       ]>�@���`�?��;Cb���yb!�sP��`�@�f����C��|�e������B��Ab�9�#*�B��8@i��C�C�i�B�����'@�-����\��g3���B�3t��$�Á��A�%���#�cCAs�B����#�Aq�B2ƑA7�C=��B�w�@�$�C���A�� ���W����`��苋A� �F�@�R��C��IN@Ag@�B�U��+CQ�\A�ׇ�|8���RB�y_Aȡ�²�$B��@h��A��A�](����5A�U@�p����B����1C=�*A����vA(e,z�������¥0_���A_�N�,�g�c�A&~��5��@
��>�Fg�@&��2�U�����]L       
categories[$l#L                                          	   
                                                 L       categories_nodes[$l#L                                   0   3   6L       categories_segments[$L#L                                                                                     L       categories_sizes[$L#L                                                                                    L       default_left[$U#L       ]                                                                               L       idi(L       left_children[$l#L       ]               	            ����                        !   #   %   '   )   +   -   /   1   3����   5   7   9   ;   =   ?   A   C   E����������������   G   I   K   M   O   Q   S   U����   W   Y��������   [��������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       ]H�O'Ij��IzH��
I�;ICM�I�h!Ira�I%��    H�I5�H%|hIXHx)�I�^�I�@�IQ�I�xD߿�G� I��NIW�aHV�hG+(F��CG�     F��I��I��AI�CJ)��I�IQI�7�I�K�                H�g�I��OI"�I��;H%0G�szE0�E�    A�Z�F|(         D3�                                                                                                                                                        L       parents[$l#L       ]���                                                           
   
                                                                                                                                   !   !   "   "   #   #   $   $   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   2   2   3   3   6   6L       right_children[$l#L       ]               
            ����                         "   $   &   (   *   ,   .   0   2   4����   6   8   :   <   >   @   B   D   F����������������   H   J   L   N   P   R   T   V����   X   Z��������   \��������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       ]?�V?�x�B�  >I�      ?�M�D�� >����D�� >1&�?e�D�` ?�^5=B�33   D�� @�  @      @߮   >�|�   @�ƨB�3t   >׍P>>v�B��=   >A�7>���@�p�@���B2ƑA7�C=��B�w�=�x�D�� >]/@�m>aG�@�  B     �F�@@     �IN@Ag@   ��+CQ�\A�ׇ�|8���RB�y_Aȡ�²�$B��@h��A��A�](����5A�U@�p����B����1C=�*A����vA(e,z�������¥0_���A_�N�,�g�c�A&~��5��@
��>�Fg�@&��2�U�����]L       split_indices[$l#L       ]   
   
                                                                                            	                                               
                                                                                                                                                                                          L       
split_type[$U#L       ]                                                                                  L       sum_hessian[$d#L       ]E�8 E�H D� E˸ A�  D� A�  D�  E�� @   A�  C�  B0  A`  @�  D   D(@ B�  E�� A   A   B�  C�  B  A  @�  A   ?�  @�  A�  D� D� B�  A�  B�  E*P E@ @�  ?�  @@  @�  B\  A�  Cw  C  A�  A   @   @�  @   @   A   @   @@  @   A�  ?�  Cy  C�� D  A0  A�  BT  A�  A0  B�  A   E C�  E@ C�  @�  BH  @�  A�  A�  CZ  B(  B�  A   A�  @@  @�  ?�  ?�  @�  ?�  ?�  ?�  ?�  @�  ?�  ?�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       93L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       [>
�u@  	���g?�/C1�����{�@z������
c�C�	 C?ڼ�%PECk���*�ܽ��B./��s�B��U6B3_�lCي��0xLÒs��j��C2�hÀ����(�sE@A�>�A�\Cq���~��Ñ��C���l�AjK�7cD
ְC��0P­�Bó@á�<B�bV�������`��/�CSl�E��A�?�wB
�A^�d��3<�  B���?Y�l�$B9�_������BVt�C��BO�u���A4����k������}�B�&�C4�)�`��B���d�Ak�BBc]��MAq-��ӧB+�@@Qg�@�!�m�
�S�\�m��]A��C�����L       
categories[$l#L       &                         
                            	   
                                               	   
            L       categories_nodes[$l#L                $   %   (   +   -   .L       categories_segments[$L#L                             	                                   %L       categories_sizes[$L#L                                                               L       default_left[$U#L       [                                                                               L       idi)L       left_children[$l#L       [               	                  ����                  !   #   %��������   '   )   +   -����   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K����   M   O   Q   S   U����   W   Y����������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       [H�0�IżI�V�H奡I�NkI��SI�Ib}I���G�:IG�    Inv�IR��I�?I%CJe�JU�gJXG�j?        H�ʨH�S�H�ˠG�*�    Gr�PIGSInr�I��PI�V JI�IČ�J �IO�kF�w
Gd�,G� H ��Hgؕ    F�9SH�̠F�,�E��F��    I
��I<                                                                                                                                                                L       parents[$l#L       [���                                                           	   	   
   
                                                                                                                 !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   +   +   ,   ,   -   -   .   .   /   /   1   1   2   2L       right_children[$l#L       [               
                  ����                   "   $   &��������   (   *   ,   .����   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L����   N   P   R   T   V����   X   Z����������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       [?G�>�p�>�bN?�>�  =o>ٙ�>���@�RA0  B*  C?ڼ   ?�n�>�Z?M�B�     @"�@�  B3_�l@Å@?
==��>R�C2�hBV  B�  >�A�@�  D�� >r�!A   B7��B�        >�dZ?�
=   >+­�   =�o      @�Q���`�@�  D�  �E��A�?�wB
�A^�d��3<�  B���?Y�l�$B9�_������BVt�C��BO�u���A4����k������}�B�&�C4�)�`��B���d�Ak�BBc]��MAq-��ӧB+�@@Qg�@�!�m�
�S�\�m��]A��C�����L       split_indices[$l#L       [         
            
                          
   	                                 	                      
                    
                                                                                                                                                                                                         L       
split_type[$U#L       [                                                                                   L       sum_hessian[$d#L       [E�8 E�  DH� E� B  B�  D8� E�� Cր A�  A�  ?�  B|  A  D6� E�� D� C�  B�  A`  @   @   Ap  B  A�  @�  @@  A   D4� E�p D@ C� B�  C�  BX  A�  B�  @�  @�  A   @�  A�  @@  @   A�  @�  @   @�  @   D2  A   E�� B�  C�� B�  C�  C'  A�  B\  Cu  B  Ap  B  A�  @�  A�  BX  @�  ?�  @@  @�  @   A   @   @@  @�  A�  ?�  ?�  @   A�  @   @   ?�  ?�  @�  ?�  C�  Cr  @�  @�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       91L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       ->>2�>�~��k��>NC>E�¥(���Z�@�����ć���kC�UD?�` B9��W�)>�C�A�Q���F�BQ�C6�A\�!����C��Ctn���C@|��'����ABm?:�A�[�b�����@Y�v��B����[<}@�r�C�?�,p���ƁCD%�A�U���oD@1#L       
categories[$l#L                                          	   
   L       categories_nodes[$l#L                L       categories_segments[$L#L                             L       categories_sizes[$L#L                            L       default_left[$U#L       -                                         L       idi*L       left_children[$l#L       -               	��������                        ����   ��������         !   #   %   '   )   +������������������������������������������������������������������������L       loss_changes[$d#L       -H�eH���EހH�nI a�        I.�I�͠GbղF��`I���I��_I��pI���    E��        I���I��IK��J#��J3:WI�	$JYvI�s                                                                        L       parents[$l#L       -���                                               	   	   
   
                                                                              L       right_children[$l#L       -               
��������                        ����   ��������          "   $   &   (   *   ,������������������������������������������������������������������������L       split_conditions[$d#L       -CD  C4     >���>�V¥(���Z�>��7=ě�B�  B
ffB�  Bb  @�  =���A�Q�   BQ�C6�B�  B�  A��   @�  >R�>�v�>����ABm?:�A�[�b�����@Y�v��B����[<}@�r�C�?�,p���ƁCD%�A�U���oD@1#L       split_indices[$l#L       -               
                                                                  	                                                                              L       
split_type[$U#L       -                                          L       sum_hessian[$d#L       -E�8 E� @�  E�� A   @@  @   E�x E6� @�  @@  Ej� C�� CЀ E� @@  @   ?�  @   EI  D� Cu  C  A�  C�  B  EP ?�  ?�  E;� CR  B4  C�� Cf  Ap  B�  BP  A`  @@  C  C�  @�  A�  C�� E� L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       45L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       }>E��BI�@��A�����g�@�FA��aABE�B���w4��>"�DdAd�16B]�@�KC��7B�C�Z� �h��g�@�؍�mM��R��G�A�o��Q�������A���B�wBF%��S@ D ���+�LCvfB}�UC�*B����zZ�¢3n�Vu�By��/����iA�����A΀��q�C��B@(S���B�o4¡ 1��Ó{���W�Cb��B�4�O�@�S�Cx�@ڤaB��s�/t'¾_�B���A��C{�@�������p�A_o"C![#�3��Bi��C��A�/~��nA�bnA'�)���}��-�?^�?�сB�T��tp��>����9¬qB�Z¬� �������V�D}�A�	s�J�´�$C�d$B3eA!$�Bkh@��C^A�0�B�v1A\���{���w��:&��W��!g@4ʣ�(�C&�[A<9�A2���aZ�B#����Aj����B�X����gL       
categories[$l#L       +                                                                        	   
                                                  	   
      L       categories_nodes[$l#L       	   	            !   "   )   .   >L       categories_segments[$L#L       	                                                                !L       categories_sizes[$L#L       	                                                               
L       default_left[$U#L       }                                                                                                             L       idi+L       left_children[$l#L       }               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K����   M   O   Q   S   U   W   Y   [   ]   _   a   c   e   g   i   k   m   o   q   s   u   w   y   {��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       }H�d�I��fI'��I7!�I&Z�I�!I���I@]<JdI�{I��IN� I��I9�tIo�HIMH�H���I�vJ1�I��I.I���I�#rIJzxJ+lI��kI��IEe
IF�bI��dIi0�I��I��G�w�I?XI<9�I�>�H�H�    I��$IqmH�d�I��J��IN��H�K�IK�I���I�yI��OI�<�I�a�I�HԹIj�H��mH`�I�EIN,IrC>I��PI\?I�&X                                                                                                                                                                                                                                                        L       parents[$l#L       }���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   $   $   %   %   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <   =   =   >   >L       right_children[$l#L       }               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L����   N   P   R   T   V   X   Z   \   ^   `   b   d   f   h   j   l   n   p   r   t   v   x   z   |��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       }A  D�@ D�� B��=?p�?�B
ffD�� @�     ?�VB�     >T��>ؓu?�A�@�  ?�n�   >�?}B[��@   B�  ?o\)A�  >���>�P   @�=q>�7LB0  Bl  Bt        ?;d@@  B�  C�*@   @�m   @��R?���D�� @�     ?C�
@@  >�Q�@�  B�  ?��>:^5B�  @E�A  @�\)@�z�A��>�E�>�9X   @ڤaB��s�/t'¾_�B���A��C{�@�������p�A_o"C![#�3��Bi��C��A�/~��nA�bnA'�)���}��-�?^�?�сB�T��tp��>����9¬qB�Z¬� �������V�D}�A�	s�J�´�$C�d$B3eA!$�Bkh@��C^A�0�B�v1A\���{���w��:&��W��!g@4ʣ�(�C&�[A<9�A2���aZ�B#����Aj����B�X����gL       split_indices[$l#L       }                  
                
                            	                  	                                                
         
                   	         	   	                     
                                                                                                                                                                                                                                                               L       
split_type[$U#L       }                                                                                                                    L       sum_hessian[$d#L       }E�8 DՀ E�� D	� D�� Ep@ D�� C�  B�  C�  D3  E� D�� C�  D�  C� @�  B�  A`  C_  C[  D � CI  D�  C�  D�� Cx  B�  C.  D�� C;  Cf  Ci  @@  @�  A�  B(  A   @�  B�  C  C&  BT  CX  C�� C+  A�  D�� D$� C�  A   DP@ C�� B  CQ  B�  A�  C!  AP  D  BH  B�  B�  CK  A�  CV  A�  @   ?�  @   @   A  Ap  B  A   @@  @�  ?�  B�  B�  A�  A�  C  A�  A�  C'  BD  @�  C�� C%  @�  @�  A�  D�@ CK  Ca  C�  C�  B   @@  @�  D>  B�  C  B�  A0  A�  C6  A�  B@  A�  A�  @   B�  B  @�  A  Dz@ A�  A`  B  B`  A   B�  B  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       125L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       y>kH�A��࿟��B�R���<J4<̴o@���Cb��A�f���A����)j;Cߞ�t
;��]B҄#C���Bz5l�Lp�Bg���2�D��B�s��lø.,�@'�D%��?�Q�yLXC��p�C������CY3D6@��%ׄC�ӶB�vdóu�C��?���B��`��C{�c��C:�ZV�CF�!�VФ�+��#.C/���<��S�CLvHD:�B��H�>���ϻB-���`�C�����Bc���V��?$V4B屨A�)�²vdBb� �B�P�C�7�¥��B�lD�-�wB�FB���G��D�a�i@��p�B{�[�,	�A�B#Y�̩B�W�§-��!usB���B�К�'�¬��B��@�2�AP64���g��^C@�:A�T�ªh�B4JtµU�A޵��c��C �Cz�HA���B�yB���¿��B	�Y°���c<��{B$��������eL       
categories[$l#L              	               L       categories_nodes[$l#L          
            +L       categories_segments[$L#L                                           L       categories_sizes[$L#L                                          L       default_left[$U#L       y                                                                                                                 L       idi,L       left_children[$l#L       y               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y��������   [   ]����   _   a   c   e   g   i   k   m   o   q   s   u   w����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       yHi�cI���I/tI�_�I�r�I�y�I[v�I{]yI���I�RqI�;�I88�Iz��J"�"IVUmI;��In�UJFdI��I�0qIW+�I�IQ�IW?pI���H�ӀI�I���IbI��H��JH�}�I1'I(�>IN_<H��{I}3I���IB7�I�zI!��IX�~IB�+H��I��        I�0)I��    IJ$Gc�Hc+�H��uIn�I6�:I���H�0H��IK�H�I�eI��                                                                                                                                                                                                                                        L       parents[$l#L       y���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   /   /   0   0   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <   =   =   >   >L       right_children[$l#L       y               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X   Z��������   \   ^����   `   b   d   f   h   j   l   n   p   r   t   v   x����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       yD�` >-VD�� >$�@@  @  D�` BM�>��=��
   B�  =�>�$�D� =�9X=��>�"�=�Q�?�z�>���B(G�   @�  =��   >+BL  >>v�>I�D�`    ?:�H<���>��>��?�{?S�>C�D�` B.  @@  >aG�   <uC{�c��=�
==q��CF�!B�  =��m=ix�=��@�  @�G�=���@�  B'
=>2-B  ?+C�D�� C�����Bc���V��?$V4B屨A�)�²vdBb� �B�P�C�7�¥��B�lD�-�wB�FB���G��D�a�i@��p�B{�[�,	�A�B#Y�̩B�W�§-��!usB���B�К�'�¬��B��@�2�AP64���g��^C@�:A�T�ªh�B4JtµU�A޵��c��C �Cz�HA���B�yB���¿��B	�Y°���c<��{B$��������eL       split_indices[$l#L       y      	      	                                          
         
                                                
      
   	            	                                                       
                                                                                                                                                                                                                                                 L       
split_type[$U#L       y                                                                                                                    L       sum_hessian[$d#L       yE�8 Cր E�� C  C�  C   E�� B�  B�  C;  B�  B�  Bd  B0  E�p B4  B@  A�  B  A�  C"  B�  @@  BL  A�  A�  B   B  A   A�  Eɸ @@  B(  A�  A�  A�  AP  A�  A�  A   A�  Bp  B�  A�  Bl  @   ?�  A�  A�  ?�  A�  @�  A@  A@  A�  A�  Ap  @�  @@  A�  @�  C6  E� @   ?�  @�  B  @�  A`  A�  @�  A�  ?�  @�  A   Ap  @@  @@  Ap  @�  @�  @�  A@  A0  BD  A�  B�  Ap  @�  @�  BT  A   A�  @   A�  A�  @   @@  @   ?�  A0  ?�  A0  A�  @�  A@  @�  A  @�  @�  ?�  ?�  @   @�  A0  @�  @   B�  B�  @@  E�� L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       121L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       E>���?&��¥�*>��B�l�B66ÓB�?nΛ��A��C�D{��Czp��#-��)�ºk~?�{�����h	�C#��v�CLZ�B��xC��x��\D�1Md�Q���&��C��-A`�7���~B�����I�Ñ�1�6� Bh΃���4B�	£U�A��?�94Bԁ$A�,m�:����c��9�£ӰA��C�����AZc�ʠ�������jA����B��B?�c��-��ˤA�
��1v*A��M@����9��z\¸^0�~V���Aę�L       
categories[$l#L                                                         	   
                L       categories_nodes[$l#L                         "   %   &L       categories_segments[$L#L                                                                L       categories_sizes[$L#L                                                               L       default_left[$U#L       E                                                         L       idi-L       left_children[$l#L       E               	                     ����   ����            !   #   %����   '   )   +��������   -   /   1   3   5   7   9   ;��������   =   ?����������������   A   C������������������������������������������������������������������������������������������������L       loss_changes[$d#L       EHKzH^��I=��H���I# zI)T!G�y�H�c:H���H$
H�@~H�
�    FBu�    IcȿHQ��H�7bH/�G6B0Gw�>    E�r`F�T(H )�        H���H�dI��
H�H1"XHy7�H� Gz;!        D�>�FH�0                G�LG��!                                                                                                L       parents[$l#L       E���                                                           	   	   
   
                                                                                                           !   !   "   "   %   %   &   &   +   +   ,   ,L       right_children[$l#L       E               
                     ����   ����             "   $   &����   (   *   ,��������   .   0   2   4   6   8   :   <��������   >   @����������������   B   D������������������������������������������������������������������������������������������������L       split_conditions[$d#L       E@��\@�v�?	��@���A��BT     <���   >�+B2  =��Czp@@  ��)�>���>;dZ?��      @�  CLZ�@@     =�h�1Md�Q��?��HB33?7K�>�33@   @�  A0     Bh΃���4      A��?�94Bԁ$A�,mAQ�A����9�£ӰA��C�����AZc�ʠ�������jA����B��B?�c��-��ˤA�
��1v*A��M@����9��z\¸^0�~V���Aę�L       split_indices[$l#L       E                               	      	                                                                                                                                                                                                                L       
split_type[$U#L       E                                                             L       sum_hessian[$d#L       EE�8 E�P A�  E�x A�  A�  A   Eٸ B`  A�  @�  A�  @   @�  @�  A�  E�� B,  AP  @�  A�  @   @@  @   Ap  @@  ?�  A�  @�  D�� E�� A�  A�  A   @@  @�  ?�  @�  A0  @   ?�  ?�  ?�  @�  A   A0  A`  @   @   D� D  B�  E�� @@  A�  A�  @   @�  @�  @   ?�  ?�  @�  @�  @�  @@  @�  @�  @�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       69L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       u>i.@ކ����}�Qg�A������"��c�A�� A��eCS�AB�i
�		�Aq ��L�wA����&��C�
�A��'¤�B�SC�kB6\BV�SD;(B�&��?ՓA\�DGc��i��u Bp�����F��Ë������C�B	�� N��z�U FB�\=�0��C-D)��C����d�wC���CES�BRB��+C����Z-C���A���W4Co�A�g��A��C��\���_0���DB:A!�d��c,��5�����D�h�'�BE��C9��B?��@������}���E>�G��c;������3&@Z��B%�����A�'�C���}$�Co��AtqgB��Z���̬�Bȳ'B�w*AP�B������@`���_)�C%2*��HZ@���§�~C	��A�P���ohAT�����"CP�� ��ҏ�B�%B�Th�����p?�/�L       
categories[$l#L                         
                           
                          	          L       categories_nodes[$l#L       	      	                   $   =L       categories_segments[$L#L       	                      	       
                                   L       categories_sizes[$L#L       	                                                               L       default_left[$U#L       u                                                                                                L       idi.L       left_children[$l#L       u               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E����   G   I   K   M   O   Q   S   U   W   Y   [   ]   _��������   a   c   e   g   i   k��������   m   o   q   s������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       uH��JIaBI+��I)�I��I��&I#�I���I�(9I˭�I��Iw�I�� Ik%(INZ�I���I�U|I�Ib'TIKXJ��IϴI�d1H�� Fr�Io�I��DI)��H��"I�n�J�jI��I�[I�/�I�p    H���I�P>I�`�I
�Ija�I�7�IƂ+IDV"IS� IZ�|I��H��eH�        G��I���I�T�G�{�I=��IZ�        I�sRJ��I�s�H�@�                                                                                                                                                                                                                        L       parents[$l#L       u���                                                           	   	   
   
                                                                                                                                         !   !   "   "   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   3   3   4   4   5   5   6   6   7   7   8   8   ;   ;   <   <   =   =   >   >L       right_children[$l#L       u               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F����   H   J   L   N   P   R   T   V   X   Z   \   ^   `��������   b   d   f   h   j   l��������   n   p   r   t������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       u?WK�?%�?bJ>uB�     D�� ?�(�=�o   >�$�Bt  B�\B�  B  @@  >k�?��HB  Bd  >�
=>Z�D�     B�     A        A�  ?�^=�S�   B�  B�  ����   >�=q?�A   >I�^@�  >��!D�  @�  ? �A0  D�` =���CES�BRB@@  >�+>�>��>�?}D�  Co�A�g�D�� >��   >��u���DB:A!�d��c,��5�����D�h�'�BE��C9��B?��@������}���E>�G��c;������3&@Z��B%�����A�'�C���}$�Co��AtqgB��Z���̬�Bȳ'B�w*AP�B������@`���_)�C%2*��HZ@���§�~C	��A�P���ohAT�����"CP�� ��ҏ�B�%B�Th�����p?�/�L       split_indices[$l#L       u                                                                                                                      
                                 	                 	                       	      	                                                                                                                                                                                                                        L       
split_type[$U#L       u                                                                                                            L       sum_hessian[$d#L       uE�8 EI� Ep� E� DF� C$  Ef� D�� Dj� D8� B\  B<  B�  D�� E� D-  DH  A  Dh@ C	  D� A�  A�  B0  @@  A�  B�  D�� @   E� B�  C�  C�  DB� A�  @   @�  D2  CY  B�  B  CȀ CI  Ap  A0  Ap  A`  A�  A�  @   ?�  A@  A0  B�  @�  D�� C  ?�  ?�  E� B,  B�  A   C  CM  C4  C,  D@� A  A�  @�  @@  @�  B�  D@ CO  A   B�  A�  AP  A�  C3  C^  B�  B�  @�  A   A  @   A0  @�  A@  @   A   Ap  @@  A�  @�  @�  @�  @�  A�  B�  @   @   D
@ D'  C  @   B�  E` A�  A�  @�  B�  @�  @�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       117L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       m>���?���p���B��B��Y֞��FBs��B^�ã�AsC�zÈ�~� �*?J���B,@C)b>���B��&B.���h���CWOTD���98 ���Af�9C)(�eeH����B��7�>�AuiC���
�ä��BWb�V3,C~��Cl���P|@äA���8�B���Az�Bْ���? C@za@dgB�R�s��o+ ��B՝��wCi�u��.��-��.Q�����.��hpB��Bo���d'�B�p���;�?��B���A�EI�|����&������ZB|4lA�h�;$C 0)@�H�B��mA��A�/Z�̧��4AnݚA�h������Z��Z�AYS�����BvJz@�����g@���A/]4�]!B5_���tB�7FA��4?Ջ4��4��B�M�A:���Fs�L       
categories[$l#L                                             	   
                          L       categories_nodes[$l#L          ,   0   3   5   6   7   :L       categories_segments[$L#L                                                         L       categories_sizes[$L#L                                                        L       default_left[$U#L       m                                                                                                L       idi/L       left_children[$l#L       m               	                                    !   #����   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S����   U   W   Y����   [��������   ]����   _   a   c����   e   g   i   k������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       mHY�pH�8JIFhH�d�J��I�ISAH�~eIAS�I�� I�v�H�IC�I�v1H���I��\Iڭ"I��    J#�J@�WH��J��H��H���H�/@HgXI#sxHHa�G��hH�O�Il��J7�,I���I�N^I�I>�$IO|(J�J;�J>U�G�H<��    F���G��`HYPD    FJ�F        G20Z    F`f�I|�G��?    FJ�`D��:IA�I1                                                                                                                                                                                                L       parents[$l#L       m���                                                           	   	   
   
                                                                                                                                   !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   ,   ,   -   -   .   .   0   0   3   3   5   5   6   6   7   7   9   9   :   :   ;   ;   <   <L       right_children[$l#L       m               
                                     "   $����   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T����   V   X   Z����   \��������   ^����   `   b   d����   f   h   j   l������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       m@�  B�=q>\)A@  A  >�M�>8Q�B�  B�  A�  D�� D�� D�� B�  >j~�B�  >I�>)��C)b>@w�>ix�>H�9D�  >:^5A   A   D�@ >C�@�  C  >W
=B�  >���=�;d>L��>o@@  @@  @   >9XB  A`  B̊=äA�   >��>C��Bْ�   C@za@dg   s�         �w@�     A0  @�  ����.��hpB��Bo���d'�B�p���;�?��B���A�EI�|����&������ZB|4lA�h�;$C 0)@�H�B��mA��A�/Z�̧��4AnݚA�h������Z��Z�AYS�����BvJz@�����g@���A/]4�]!B5_���tB�7FA��4?Ջ4��4��B�M�A:���Fs�L       split_indices[$l#L       m                  	                                                       	            	         	                                              
   	                                                                                                                                                                                                                                                   L       
split_type[$U#L       m                                                                                                      L       sum_hessian[$d#L       mE�8 E�P C  E�� C�  B  B�  E̘ B�  C�� Ap  A�  A   A�  B�  E�h C�  B�  @   B�  C1  @�  A   A�  @�  @�  @�  A   A   @�  B�  E�� B�  B�  Cc  A�  B$  A�  B�  B�  B�  @�  @@  @�  @�  A@  A  @�  @@  @�  ?�  @�  ?�  @@  @�  @�  @   @�  @   A�  B�  E�X B4  B  BP  A0  B�  B  C@  A�  A`  A�  Ap  A   A`  B0  B0  B�  A�  B0  B  @@  ?�  ?�  @   @   @   A   @�  ?�  A   ?�  @   ?�  @@  @   ?�  ?�  @�  @�  ?�  @�  ?�  ?�  ?�  A�  @@  BP  A�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       109L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       s>0	~A����e���6�B������Y{�f�B��MB+\OC;�3É�@��#Co]��c��B���C.���!V�A�9@Cf��DBo9B���C�@���-�Ñ4B4$�C����)WuB{��2lAW����en��״�|�C�d>��3C<OÜ�AB�vI�欯B�ӓD,�DqZ:C![��:ZB�b.A����X������[�B\��H2tB�V�B��kD-�c�«��B�ʟ�Ѽ��&-������B�A�A��O�3�)�C�B�G��2�NBp�@Ě�B/����vA~]B�ۍ��fXB��
PB9�BCd�zBH�MC�EfB�R��r/B�L��o �5�B �W���0��J��	�M��kMB���>��@�k��y5C�iA�}IB�����Cb�+Bn�'��m��ـ�hn�A���]�ZA�ʓA΋��ȑ�(���_L       
categories[$l#L       2                         	                                                    	   
                        	                                      	   
         L       categories_nodes[$l#L                               %   +   1   3   4   8L       categories_segments[$L#L                                                                                     "       #       $L       categories_sizes[$L#L                                                                                                  L       default_left[$U#L       s                                                                                               L       idi0L       left_children[$l#L       s               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A��������   C   E   G   I   K   M   O   Q   S����   U   W��������   Y   [   ]   _   a   c   e   g����   i   k   m   o   q����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       sH���I�G0I
��I���I_9I��I3�I]qI��I��JF��J��IA��I�D�H���InB�G���JN I��{IF-I��II�rIx#jF��I��H��PIDcI���G!�IF}6H�'~I�
I��J        I��H��nF�WxI��I�#I"HڻPG���E�`     I�^�H��Z        HW/�I�(G��F��I(��I5.H�FxHhw�    E>ߐI+ƫI��IT��H�8/                                                                                                                                                                                                                L       parents[$l#L       s���                                                           	   	   
   
                                                                                                                                         #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   -   -   .   .   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   :   :   ;   ;   <   <   =   =   >   >L       right_children[$l#L       s               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B��������   D   F   H   J   L   N   P   R   T����   V   X��������   Z   \   ^   `   b   d   f   h����   j   l   n   p   r����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       s=�t�>��\=��
?�B��{D�� =��>��7@�  >\B�     >t�   >�->T��   ?.�?�   Ap  @�  D�        A  ?�=q   >���@_\)>o��=��B
ff��״�|�D�  =�P   =���?�@�?��A      :D�� @�  B�b.A���   D�`       =��PD�� @�     c�D�� B  @�  D�@ >�  �B�A�A��O�3�)�C�B�G��2�NBp�@Ě�B/����vA~]B�ۍ��fXB��
PB9�BCd�zBH�MC�EfB�R��r/B�L��o �5�B �W���0��J��	�M��kMB���>��@�k��y5C�iA�}IB�����Cb�+Bn�'��m��ـ�hn�A���]�ZA�ʓA΋��ȑ�(���_L       split_indices[$l#L       s      	      
            	               
                                                    
                                 	                                                                                                                                                                                                                                                                                              L       
split_type[$U#L       s                                                                                                      L       sum_hessian[$d#L       sE�8 D� Eɠ C�  C�� B�  E�� C�� B�  Cd  BT  A�  B�  A�  E�� C�  @�  B|  A�  CJ  A�  @�  B8  @�  A�  @�  Bh  A�  A   CU  E�8 C   C  ?�  @�  A�  B  @�  A`  B�  B�  A�  @�  @�  ?�  B  A   @@  ?�  A  A`  @�  @   A   B@  A`  @�  @@  @�  C5  B   C�� E�  B   B�  A�  B�  @@  A�  @@  A�  @�  ?�  @   A@  B�  @�  B�  A�  @@  A�  @�  ?�  @�  ?�  A   A�  A   @   @�  @�  @   A@  @�  ?�  ?�  ?�  @�  @�  @@  B4  @�  @�  @�  @   @�  ?�  B$  C  A�  A  B�  C   A�  E�` L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       115L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       s>@��@����Y@���������4x���f@��C���q2SÄ���D+�Â532?�!A���fVC`O\Ï�A��ҍ�F���=M?�T+�C �u@�����DDA���x��e��B��;�Ɋ�A�C�N��A䉣C����,�C�j��j�CĬzb�Xʘ�vh�Ì�O¶�hC	�s¯ZmCmB�`$p�69�'���%e�B�r��5�V�*C����B6�3C���?T*x��
]B 0@]�U��p�'lbA?q��Sc�Ѹ�C�B�����^Ai C9���n�uA�B�9�A�'�XWEA����z�k��� I�u��2:@º���g � ��8��Bn� �AuY��3Y�B�P��(���[��t�B�mX¤i�Ì9������E	B�����d�Bo!����<�\�����?���C.y���U@^D�B����CrL�BJ�L       
categories[$l#L                                      	   
                                              	   
                 L       categories_nodes[$l#L                             %   *L       categories_segments[$L#L                                                                L       categories_sizes[$L#L                                                               L       default_left[$U#L       s                                                                                                       L       idi1L       left_children[$l#L       s               	                                    !   #   %   '   )   +����   -����   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c   e   g   i   k   m   o   q��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       sHl��IT��I��5I['8H��HI���IB��H���J�VHs��H��xIO��I�`�I�@�I;�IT�hI�b�I�Q�I�Hv2G��G҂�    H��f    IO�J�I�0FIv��IS�1IbY�IA1UI��*I��CI7I|I���H��rH,��IׄHKoHGlsG2pFAPG5'F��\G|BHHo�bH���GoʀI��I���I ��Iv�9H��I�(\J}�IL�XI<��IXv�                                                                                                                                                                                                                                L       parents[$l#L       s���                                                           	   	   
   
                                                                                                                             !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   :   :L       right_children[$l#L       s               
                                     "   $   &   (   *   ,����   .����   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d   f   h   j   l   n   p   r��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       s@�Q�@BM�@��H@�{?o\)   > Ĝ>���B�  @�  @�  B�33B4(�D�  A0  ?��?ƨ   >+   >��@@  �=M?@@  C �u@      =�h   >49X@[o?��   Bh  B�  =�\)D��    B�  @   @_�wA��H   > Ĝ?K�A�  ?�jA�  @   A�  >7K�=��?#�
?�B;��@�?�%@�{=��?T*x��
]B 0@]�U��p�'lbA?q��Sc�Ѹ�C�B�����^Ai C9���n�uA�B�9�A�'�XWEA����z�k��� I�u��2:@º���g � ��8��Bn� �AuY��3Y�B�P��(���[��t�B�mX¤i�Ì9������E	B�����d�Bo!����<�\�����?���C.y���U@^D�B����CrL�BJ�L       split_indices[$l#L       s               
                                  
          	      
                                                                                                   
                  	                                                                                                                                                                                                                                L       
split_type[$U#L       s                                                                                                           L       sum_hessian[$d#L       sE�8 E� E@ E�� BH  B�  E@ E�� BT  B  Ap  B4  B  CB  D�@ Ev0 DF@ B0  A  A�  A`  A`  ?�  B(  @@  A`  A�  B�  B�  D� C  E%� D�` C� C�  A�  A�  @   @�  A   AP  A   @�  @�  @�  @�  B  @�  @�  A   AP  A�  Bl  BP  B|  B,  D�@ C   AP  E� C  Cp  D�` C�� B�  C�  A�  @   A�  @@  A`  ?�  ?�  @@  @�  @   @�  @�  @�  ?�  @�  @@  @@  ?�  @�  @@  @�  @   @�  A�  A  ?�  @�  @�  @@  @�  @@  @�  @�  Ap  @�  A�  A�  @�  B<  A�  B  B  A  D=@ D�� Bp  B�  @   A0  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       115L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       /=�uY>�CX�-G=�yBCb���9N��8UA2�7� .�B��B���T���Q g@u���@*��p�A�-���>��@�gB�d��ێ���,��c'BtHF@�@��$��;FAc�����B�����k�A����7YAw��C�d��g�AZ�AHO��a���EF���@��}��V����p�^L       
categories[$l#L                                             	         L       categories_nodes[$l#L                L       categories_segments[$L#L                             L       categories_sizes[$L#L                            L       default_left[$U#L       /                                             L       idi2L       left_children[$l#L       /               	            ����      ������������            ����������������      !   #   %   '   )   +   -����������������������������������������������������������������L       loss_changes[$d#L       /HF�bH�+�G�HEǦG���F�� E�I��I��    E�:HD�             I~�I5<VI���H���                H�>I�*XI��`I��I�VoJ~I���J��                                                                L       parents[$l#L       /���                                                           
   
                                                                              L       right_children[$l#L       /               
            ����      ������������            ����������������       "   $   &   (   *   ,   .����������������������������������������������������������������L       split_conditions[$d#L       /CB  C4  =t�?���D�@    B�  >�P?�G�B��B  D�@ �Q g@u���@*�      D�  >R�@�gB�d��ێ��=>�+?E�Bb  ?:^5B4  @�  B0  B�����k�A����7YAw��C�d��g�AZ�AHO��a���EF���@��}��V����p�^L       split_indices[$l#L       /                                                               	                         
                                                                               L       
split_type[$U#L       /                                            L       sum_hessian[$d#L       /E�8 E�� A   E�� @�  @�  @   D�� E�0 ?�  @�  @�  ?�  ?�  ?�  Cm  D�� Cހ E�H ?�  @@  @   @@  CA  B0  C�� DA  C�  C  D�  Ev� @�  C=  A�  A�  C�� @�  D� Cn  CI  B�  B�  A�  D�  B�  Es  BX  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       47L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       s=S�9@D6�N����FZA�a�«s��I�UA�� O���hBu���B����MC�)��gB �	�;���TAiz����K�7`gBݠ��Y��B0!#BE�CLT"�w��B�U�f[C���A����ES'B��@��wÎ�B��WBCzN�Jx�A�H4�c�4�#êEA�A�B��(����C1ҕ�(��Ñ�B�T�zVCxS��R��B����jDX�B �)AX�UD����[A����M.x����A�΍�F�@�ܤ�*����O�B���D�B8�R�D,��ѿ�xA����Ң�+&±������d�Ø���QB"�p����B���@���"�BL}�A���B�`��A��B��+T �MJB$y��.�4�(�xZB��+Az�gA���\βA箈�D�g�Gu�AJ��A3�@CWg5B��;@'����tB��Cwy2Bp+ZL       
categories[$l#L                                   	                                                             L       categories_nodes[$l#L                         "   2   5   8   9   :L       categories_segments[$L#L                      
                                                               L       categories_sizes[$L#L              
                                                                      L       default_left[$U#L       s                                                                                              L       idi3L       left_children[$l#L       s               	                                    !   #   %   '   )   +   -   /   1   3����   5   7����   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c   e   g   i   k   m   o   q��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       sH1ȣH�BI"��H�կI��ZI��FI�m�I��I1�%I�2eI�b�I�j�I4M^I�I��I��;I�AI��I1eBIB��I�u�I��J�I:yHv�CI�    I"�I���    ISDI��I��\I��I�I�=�H*Q�I�:�Ik��IWrGCJ�IJ*{I�g�H��H���I�5�J��H���IT�hH<]�GBH
�HȟtI,�7I0�H�0TH���G>�qI5R�                                                                                                                                                                                                                                L       parents[$l#L       s���                                                           	   	   
   
                                                                                                                             !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   :   :L       right_children[$l#L       s               
                                     "   $   &   (   *   ,   .   0   2   4����   6   8����   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d   f   h   j   l   n   p   r��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       sA   @�  =m�h>Y�>aG�?��FB�  >�;d<#�
>333B2  A   >ڟ�@;dZD�` ?MO�      >9X   B�
=@;dA0  <�1>���   CLT">�>n�f[   ?j>�ƨ>�F   B�  ?�z�>�  >��7D�  @�  BX  >6E�>��>�X?�\D�� D�@ >�5???}   >��BM�   D�  A��         ���[A����M.x����A�΍�F�@�ܤ�*����O�B���D�B8�R�D,��ѿ�xA����Ң�+&±������d�Ø���QB"�p����B���@���"�BL}�A���B�`��A��B��+T �MJB$y��.�4�(�xZB��+Az�gA���\βA箈�D�g�Gu�AJ��A3�@CWg5B��;@'����tB��Cwy2Bp+ZL       split_indices[$l#L       s                        	                                  
                                	             
                                     	            
                                                                                                                                                                                                                                                                L       
split_type[$U#L       s                                                                                                        L       sum_hessian[$d#L       sE�8 E�� Dj� E�p DK� B�  DO@ Ep E>p C�  C�  B�  A�  DK� A`  D�� D@  A�  E= C�� B�  C1  C�� Bp  A�  A�  ?�  DB@ B  @@  A0  Dz� C�� C�  C�  A�  @�  CM  E0@ C�� A@  B�  A�  C  B  B�  C*  A�  B(  A�  @�  A  A�  B�  D+@ @�  B  @   A  DC� C[  B�  C̀ C�  A�  C�  A�  A@  @�  @@  @@  B�  B�  Cπ EP B�  CA  @�  @�  Bh  @�  @   A�  AP  C  A@  A�  B\  B  B�  B@  A   A   A�  A�  Ap  @   @   @   @�  @@  A  A   B�  A0  D  B�  ?�  @@  @   B   ?�  ?�  @�  @�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       115L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       }=� @�]�����A�O9������<]?��f�ltB��£k�@�����NO@����%D���C[AޗCi���})�CĢA��H��+�A��:���6�B5�@R�YC�F	B^��+����B��B�!�C|����Bo�C�I@��,���aBh�>áf��F�B} ��w^B����]@g��C�%BlBH�B[�]ʠ�g�uCX>��k[P��3�B��vD�B�x�CG e½%u� ����@��I�sw�Bk+@�EdB��u@C����m���gB���A¸B�YC3U��3��B��#@�2$E�>��KB�+��\'�	���#,(B\V=@;��A�V�>��p��A��-�`���y�A����_OB!��AxwCH�A�������`���b�8���B[�NB0����ҿ���C*���q-mAwg9>.���DB	��>C]
A����W�Bt9�B���zpB�QO�;_u£���4�J�~����*L       
categories[$l#L       7                    	                     	                               	   
                           
                                                        	   
          L       categories_nodes[$l#L       
       	               %   )   <   =L       categories_segments[$L#L       
                             	                     $       %       )       6L       categories_sizes[$L#L       
                                                                      L       default_left[$U#L       }                                                                                                                 L       idi4L       left_children[$l#L       }               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C����   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c   e   g   i   k   m   o   q   s   u   w   y   {��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       }H:��H� �H�zI^�rI9 Ix�H�B�I�*�Itq�I=�ICs�I�}!I�A�Ir�I0�9I��XIx�IWrI��I� I\��Ik��IǔIw�II���I�lIa��It�I���I�WI�ΘH�>H�<:    If�I7�tI�lRI4PpI�.IF��I�H�E�I���Ib@2H�rnI)��I~��J=�H˟I8lI��JYcI�&�I'=�II�+�H?�PH*r�IT�PIL�I&��H��w                                                                                                                                                                                                                                                        L       parents[$l#L       }���                                                           	   	   
   
                                                                                                                                         !   !   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <   =   =   >   >L       right_children[$l#L       }               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D����   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d   f   h   j   l   n   p   r   t   v   x   z   |��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       }   >.{>�@�  ><j=�@5�B  @�   @�Q�D�� D�� @/
=>�K�?�P>'�=<j@�  >n��?��A      =��   B~>���@�(�   D�  D��    >p��>�$�C|��>�=qD��    A@  D�� A�     @@  @�  >��? Ĝ?KC�>���B�  ?��yD�� Bd  =���BH��A�  @߮A�  B6  B33?�$�      @@  @��I�sw�Bk+@�EdB��u@C����m���gB���A¸B�YC3U��3��B��#@�2$E�>��KB�+��\'�	���#,(B\V=@;��A�V�>��p��A��-�`���y�A����_OB!��AxwCH�A�������`���b�8���B[�NB0����ҿ���C*���q-mAwg9>.���DB	��>C]
A����W�Bt9�B���zpB�QO�;_u£���4�J�~����*L       split_indices[$l#L       }                                                            	                                                     
                               	   	                                       
                                                                                                                                                                                                                                                                  L       
split_type[$U#L       }                                                                                                                   L       sum_hessian[$d#L       }E�8 EC0 Ew@ Dp� E  DM� EC� CJ  D>@ B�  E   D  C�� E5� Ce  C&  B  D-  B�  B�  B  D�  DH  C�  C6  CX  B�  E4� AP  Bd  C,  B�  B,  B  ?�  A�  D%� A�  B   B  B$  A�  A�  DZ� C�� C  D$� C�  B�  B�  B�  C  B�  A�  B(  E)� C2  @@  A   A�  A�  BD  B�  B$  B�  Ap  A�  AP  A�  A  A�  A�  D!@ A�  AP  B  @@  A�  A�  B  @�  A  AP  A   @�  D@ C�  C�  B�  B�  B4  D� C  Cg  BD  B�  AP  B\  A   B�  B  B�  A�  A�  BD  A�  A  A�  A�  E'0 B  C  A�  @   ?�  @@  @�  A�  @�  @�  A�  A�  A�  A`  B�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       125L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       Q>b�unB")� ��B���@�v�C5�:?��q��b���0Bb���C~�d����B6�G��7qB������yC M2�\�A'ɴ½�C�D�@I������)BoCM$���e��B�����C��`�&��CA���������C�.����nKB�P���D4� T�C8;DC�LAF����P ���_Brþ�4��B����I0o�<}�B;y�hK��%�B9��ĪoA�#r�I��B�Ag��B����w���PD�2l�C!�RA̰�A�5���@�� �?�&Bw����A���B���=�g��]gL       
categories[$l#L       9                             
                                           	   
                                            	   
                                   	   
                  L       categories_nodes[$l#L          	                     "   %   &   .L       categories_segments[$L#L                                                                *       +       6       7L       categories_sizes[$L#L                                                                                    L       default_left[$U#L       Q                                                              L       idi5L       left_children[$l#L       Q            ����   	                                    !   #   %   '����   )   +   -   /   1   3   5   7   9   ;   =����   ?   A   C   E   G   I   K��������   M��������   O����������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       QH6�ZHndIo�H|$f    I��H�2�H���Ir�I�I�H�_4F�zkH�p�I-�(J�]I@WI;?�H��DG�x�I8�DHXl    D�h�H^PE���I)�H�6J[i�I
��I,XI|��H�~HGu�X    H���GL��G��I$�@H��HJ�|H�!�        G�P�        C�5�                                                                                                                                        L       parents[$l#L       Q���                                                     	   	   
   
                                                                                                                                   "   "   #   #   $   $   %   %   &   &   '   '   (   (   +   +   .   .L       right_children[$l#L       Q            ����   
                                     "   $   &   (����   *   ,   .   0   2   4   6   8   :   <   >����   @   B   D   F   H   J   L��������   N��������   P����������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       Q?� �@��B�  ?�B���@@  ?ա�>�j@�Q�   ?�jD�� @�  >�^5   ?
=A`  ?�dZ@Q�7   D�� A'ɴ   @      ?���?ȴ   ?(�9B�     >A�7BH���&��   @��Bf        @��@$(���D4� T�D�� C�LAF��   ���_Brþ�4��B����I0o�<}�B;y�hK��%�B9��ĪoA�#r�I��B�Ag��B����w���PD�2l�C!�RA̰�A�5���@�� �?�&Bw����A���B���=�g��]gL       split_indices[$l#L       Q                                                        
                           	                                                                                                                                                                                                                L       
split_type[$U#L       Q                                                                      L       sum_hessian[$d#L       QE�8 Eٸ B�  E٨ @   B�  A�  Eƨ D  A�  B|  @�  A�  E�� C�  D@ B�  Ap  A@  A�  B  ?�  @�  AP  @�  E�� A�  C  Cx  C�� CJ  B�  @@  @@  A@  A  @@  AP  A@  A�  Ap  ?�  @@  A   @�  ?�  @@  E�� B  @�  A�  B�  Bt  C_  A�  C�� Bp  B�  C  A   Bh  @   ?�  A  @@  @�  @   ?�  @   @�  @�  A  @@  A0  A@  A  @�  @�  @�  ?�  @   L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       81L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       u>Gg�kGzA��B?czj��$Bwǻ�_r���tA`�;BK��A�9A���C:yV�{1Av$�86�p�B�?�A?@C2w�e̹�dsCe�C�"@8�nC������G6UBMPB�e�c�?�٦yB��PC�G���Cv�B���#B��CF��¬	�B_� ��M���N���vCo\���[B��`C�ȜB����gB�:Dۉ�
Ct5��Á>ZB�x}Z�CIA{-��wt���Y�>�s���'B	���2��EJ�C��G��5��B+&C'�hB?ɔ@��A ��zoB���@�
�B�K�A�8rA �r�ɮB �����a��8A�\��J�BF��T[�A�l��;K�B�o�Bv���'���A�g����~�����GBo��Cz<g@���B���<B��q?��ћ�9�?B4�@�B����B�@1��C�|�mχ]�L       
categories[$l#L       1                          	   
                                  	   
                          	             
                                  	   
             L       categories_nodes[$l#L             	            %   '   -L       categories_segments[$L#L                             
                            $       0L       categories_sizes[$L#L                     	                                          L       default_left[$U#L       u                                                                                                   L       idi6L       left_children[$l#L       u               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [����   ]����   _   a   c   e����   g   i   k   m����   o   q   s����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       uHTH�HzH�3.H�`�H��UI;��I+0=I+.I$%�H��H�I\�I)�4H�r�I*�H�I��I4�IE�I b:H`�IgI6��I}��H��dI�(I �H���HQ�nH��G$�PH��PI��fJ"xI�e$Ie��H8��I��I��BH��jH��)G��G�8�H̹GIP�H��N    Gے    I�aG���H��+I���    G�F0H� �HH�`G1�|    H��FH��`F��`                                                                                                                                                                                                                            L       parents[$l#L       u���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   /   /   1   1   2   2   3   3   4   4   6   6   7   7   8   8   9   9   ;   ;   <   <   =   =L       right_children[$l#L       u               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X   Z   \����   ^����   `   b   d   f����   h   j   l   n����   p   r   t����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       u?;�m?�?f$�>ě�   @�  ?�M�>���>���   B�Ǯ   Bt  ?AG�@�  >��mD�� >��   ?�>�VBh  A   @@     B:{>���B'
=B�  ?[�m@"�?.��B�  D�� @@  @�>�A�   D�     B�33@   @{@@  @�     ��[D�  C�ȜB@�?Qhs>P�`?�h�
E}  ?s33D�� D�� Z�B�\A0  A�  ��Y�>�s���'B	���2��EJ�C��G��5��B+&C'�hB?ɔ@��A ��zoB���@�
�B�K�A�8rA �r�ɮB �����a��8A�\��J�BF��T[�A�l��;K�B�o�Bv���'���A�g����~�����GBo��Cz<g@���B���<B��q?��ћ�9�?B4�@�B����B�@1��C�|�mχ]�L       split_indices[$l#L       u                                                              	                                  	                                      
                                
                                                                                                                                                                                                                                                         L       
split_type[$U#L       u                                                                                                             L       sum_hessian[$d#L       uE�8 E�� C�� Eƨ C�� C!  CH  E�� D�� Bd  C�  B�  B  B  C!  E�� B�  B�  D�@ B  A�  C�� AP  @�  B�  A�  A   A�  A0  C  A   E�� B`  A�  B�  A�  BP  D6  C�  A�  A   @�  A�  CN  B�  A0  @   @�  ?�  B�  A�  A�  A   @�  @�  A   A�  A   ?�  AP  C
  A  ?�  E�0 D� BX  @   A�  @@  Bx  A�  A�  @�  A  B,  C C�� B@  C�  A@  AP  @�  @   @�  @@  Ap  @   C=  A�  B�  A�  @   A  @@  @   A�  Bd  A�  @�  @�  A`  @�  @@  @@  ?�  @�  @�  A   A@  @�  @�  @�  A  C	  ?�  ?�  A   L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       117L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       m>Z�
�j�?�T���B0��Cݹ?G��C2��)��C X��Q+C����O�`��g@��lB�8�C���A!Hf��Bh�D'���4CgDKD��BI����i�����@f��Cs@!�����C#�C%JDBW �l1�C�`i�P��`?�B$��Cc�'�k� DR='�&��îӈ�y4B���C&�D�
�Cg��xl���"A֘����i�B�GP���KD��B���-��@�+H��"'A��B�6`A$ݮB�t�� �oA�$�C4����h�\���d�FhfBdP�����A��g�K�AB���C�b%�AM�̞l@����Y�Bz ����B���C�KBŀ�V-�ݑB
j��bx@�ό��m��'A�4N���"AO}�BŅ�u��@	��A�jC���B����MB��
��feA���CL       
categories[$l#L       	                               L       categories_nodes[$l#L                   )   3   7L       categories_segments[$L#L                                                  L       categories_sizes[$L#L                                                 L       default_left[$U#L       m                                                                                                L       idi7L       left_children[$l#L       m               	                                    !   #   %   '   )   +   -   /   1����   3   5   7   9   ;   =   ?��������   A   C   E   G   I����   K   M   O   Q��������   S   U   W   Y   [����   ]   _   a   c   e   g   i   k������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       mH4aII2�I��gI�q�I�`J �Hs`RI+��IXx�J_��H��rJ*�H��tI�I���H-O�H'/�I�^I���Iu��I��HI%��G���J8S�H��x    G��4I��I_@�I�0I>��G�/G�J�        IIŠIe8IJlII��I4��    Gk�|G]��H�G�I���        G�.LI���H�"�H��E�I�    I���I}XI���ID|J-��IG�J�7I*b�                                                                                                                                                                                                L       parents[$l#L       m���                                                           	   	   
   
                                                                                                                                   #   #   $   $   %   %   &   &   '   '   )   )   *   *   +   +   ,   ,   /   /   0   0   1   1   2   2   3   3   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <L       right_children[$l#L       m               
                                     "   $   &   (   *   ,   .   0   2����   4   6   8   :   <   >   @��������   B   D   F   H   J����   L   N   P   R��������   T   V   X   Z   \����   ^   `   b   d   f   h   j   l������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       m>2->��>9X=��
>�x�   >�t�B[��@�  B��{B�  ?�ff>t�@   >׍P>!��   B�  >%�T>��y=49XB�  @   >��>N��?��>š�@@  >��+>ؓu   D�� C%JDBW <�j@@  >���>T��>��`Cc�'   =P�`D�  >�z��y4B���>j~�>:^5@�  >u   A֘�>�A�=��   @�  >VB�  >��H@�  ��"'A��B�6`A$ݮB�t�� �oA�$�C4����h�\���d�FhfBdP�����A��g�K�AB���C�b%�AM�̞l@����Y�Bz ����B���C�KBŀ�V-�ݑB
j��bx@�ό��m��'A�4N���"AO}�BŅ�u��@	��A�jC���B����MB��
��feA���CL       split_indices[$l#L       m   
   	   
                               	                  
      
            	          
      
                                	                	              	                   	                                                                                                                                                                                                                  L       
split_type[$U#L       m                                                                                                       L       sum_hessian[$d#L       mE�8 D;@ E�� D@ C4  BL  E�8 A�  D� B�  B�  B  A@  EJ` E> A�  @�  CJ  C�  B�  A   B�  @�  A`  A�  @   A   D�@ E@ B�  E7� A  A   @�  @   C:  A�  C�� B$  B�  ?�  @   A   B�  @�  ?�  @�  A   @�  @�  A�  A   @   C�� D>@ B�  E� A   B�  A�  E6p @�  @   @�  @�  AP  C-  A0  @�  @@  C�  B  @�  A�  Bx  ?�  ?�  @   @�  A�  B`  @�  @@  @�  @   @   @�  @�  ?�  A0  A   @�  @�  C}  B0  B�  D!  Bl  A�  C�� D�` @�  @�  B�  @   @�  A�  DU  E0 L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       109L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       u>��l�P�O@� A���E2�C�S?�jS���B A9��ª�A��$C��_B���>���08C��;��-B��Ba��هv�Y��F�±G�C4�!D!0�C8}#C%ƻAK���'�@ͯ��_��\�CR��S��B)�y��8����NB�c�B��A��|���������¿���Y�A��k�,�B�{m÷p�B5�3C+.BP�C�0HC���A��+�ZIDC�Rn�2\C1�By/�6��B���>#����B	L�J��1=r�% 8B !C�Ԧ+�}�@�(�� �CK�*A��A$��BB*�A*�®�BA�m���z�+�X�>(B_^��	wo��i�µCy���BF��³|B������B�a�����m�+BJ������B�B�AE�>@B��o��A�3�C
X?�m�?T�,#�C)�@A�1M¼~A���B|���B�K��h[x?Х��f*�L       
categories[$l#L       )                   
                                                          
                                     	   
         L       categories_nodes[$l#L                      *   5   7   =L       categories_segments[$L#L                             
                                   L       categories_sizes[$L#L                     	                                          L       default_left[$U#L       u                                                                                                          L       idi8L       left_children[$l#L       u               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A��������   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _������������   a   c   e   g   i   k   m   o   q   s������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       uH0��I�$IO��I���I`��Iy��H��I�\I�#YIP��I��2I�I*�
H֥�H�LIa�Hp��Ii�I�YH��I��/H��XI]�$I�$NI�H���H*�IJ�H��ICђI�e�Hb�/I�&        I�2�I?'�I.�TI���H��TH�`�H�QH���Hɜ�I,��IC~-I��lH��%G}< H��            G�p�G�p�H[��Iy�H$�LH�.\I5��I8��I�oH���                                                                                                                                                                                                                        L       parents[$l#L       u���                                                           	   	   
   
                                                                                                                                         #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <   =   =   >   >L       right_children[$l#L       u               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B��������   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `������������   b   d   f   h   j   l   n   p   r   t������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       u=�F   =��#=\   D�� >�A�  A�  @�  ?�B   >��>A�7>��?�     @�  >�Q�?u?}B[��>�(�>�ƨ   >%@   Bt  B33>ě�D�@ >�(�D�@ @�  CR��S��?�o@�  >��>�o>�(�@@  D��    A�  ?���>t�j?��@@  @�  Bx  C+.BP�C�0H   @�     @�  @�  @�  @@  <u   Bf  ���B	L�J��1=r�% 8B !C�Ԧ+�}�@�(�� �CK�*A��A$��BB*�A*�®�BA�m���z�+�X�>(B_^��	wo��i�µCy���BF��³|B������B�a�����m�+BJ������B�B�AE�>@B��o��A�3�C
X?�m�?T�,#�C)�@A�1M¼~A���B|���B�K��h[x?Х��f*�L       split_indices[$l#L       u   	      	                                  	                   
                                                                                                                                                                                                                                                                                                                                                                 L       
split_type[$U#L       u                                                                                                             L       sum_hessian[$d#L       uE�8 D]� E�� C� CҀ B<  E� B�  C�  C  C�� A�  A�  B�  E�� B|  @�  C  C�� B�  B(  C  C  A�  A0  @�  A`  A�  BD  CՀ E�X A�  B  @@  ?�  B�  Bt  B�  C0  B�  Ap  B  A  B�  B|  B�  A�  A0  @�  A  @   @   @   A  @�  A   A�  B  A   B�  C�  B�  E�` A�  A   B   @@  A�  BP  Bd  @�  B�  @�  @�  C,  B|  B  A  @�  A�  A`  @�  @@  @�  B�  A�  B  B�  A�  A�  A   @�  @�  @@  @�  @�  @�  @�  @   @   @@  @�  @�  A   A  A�  A   ?�  A  @�  B�  A   C�  BH  B4  Eq� D�� L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       117L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       )>�)>��>�BTC)�@�� �!�c?��w���B���B���PO��=� @� ��#{��s�͔@@K��A℺? .BQ���BىA�%)¨���5H�¡�+��;�?��BrHB@��#��[������A�wA�6���/�+_?����Z?�l�L       
categories[$l#L           L       categories_nodes[$l#L          L       categories_segments[$L#L               L       categories_sizes[$L#L              L       default_left[$U#L       )                                         L       idi9L       left_children[$l#L       )               	����         ����   ��������            ��������            !   #   %����   '��������������������������������������������������������L       loss_changes[$d#L       )H-g�H&��G��HIoGB��    E���H%�eI5�    E}e�        I {�H�h�H�H��v        H�4I� �Hɝ�I���H�XYI]z    FGV�                                                        L       parents[$l#L       )���                                                     
   
                                                                  L       right_children[$l#L       )               
����         ����   ��������            ��������             "   $   &����   (��������������������������������������������������������L       split_conditions[$d#L       )CB  C4  >��7@�  D�@ @��    ?-�hB�  B���B  �PO��=� ?�B�  >�/Bճ3@K��A℺@   =C�B��{>�dZ@@  >����5H�B�  ��;�?��BrHB@��#��[������A�wA�6���/�+_?����Z?�l�L       split_indices[$l#L       )         
                
                     
                                                                                                  L       
split_type[$U#L       )                                        L       sum_hessian[$d#L       )E�8 E�� A   E�� @�  ?�  @�  E�� C  ?�  @�  @�  ?�  E�� E,  C  @�  ?�  @@  E`� D� E� Ca  B�  Bl  @   @   D%� E7� B  D  E0 A�  B�  C  B  Bd  A�  B  ?�  ?�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       41L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       u>,G�@���y@����5�pg��
n�@-�A���B���cBډ��jA_p*�G�A=>���^A��tC��CIn���_����^��P@{��B��B���:m��u��B*S��5�@שpA���L��B <�>�A����L���W��C��B���B9 B���kCB��Q�Z�uB�X�,���EZB�xA���C��Cg[ �N�*@��<��h�BPKL�<+H�1#G>(|C�� @z2�@�\�B�b$Bn[q�ʳ�B%{�;�������h>ޑ�A��dBa.��A��C�r���;B~aW��U9BFTt�,�PB��ߟB�MA�@*� #H@�DB~����N]A��2DAv�Bu��z'�A��7��l A>ۧBN	�A0k4B�*�¶2���}VA_���Z��B_B�+PA���;�!û9��������6�4��A���B��C���qo?�M�L       
categories[$l#L       0             
                                               	   
                               	   
                                                       L       categories_nodes[$l#L       
       
                &   )   6   7L       categories_segments[$L#L       
                                                  	              "       'L       categories_sizes[$L#L       
                                                                      	L       default_left[$U#L       u                                                                                                        L       idi:L       left_children[$l#L       u               	                                    !   #   %   '   )   +   -   /����   1   3   5   7   9   ;   =   ?   A   C   E����   G   I����   K   M   O   Q   S   U   W   Y   [   ]   _   a   c   e   g   i   k   m   o   q   s��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       uHXH�
H��NH��H獚I�KH��BI@��IO�zH�GHŹ�I+·IdDIT�SI	��I�I��vIp(!I���H�ԺG�SI N�I
pH��    F��H�e�IZvHI�֚I1�Ium�I�D<I�7�I��\I�� I�    H��JI�
    HKd�G��*G��VH�@�H�X|H3w\I��H��kH���F"��EH�@Gp I�ITu�Iy�eI�ɫJ@II��QI׃dI�J�IQC                                                                                                                                                                                                                                L       parents[$l#L       u���                                                           	   	   
   
                                                                                                                                   !   !   "   "   #   #   %   %   &   &   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <L       right_children[$l#L       u               
                                     "   $   &   (   *   ,   .   0����   2   4   6   8   :   <   >   @   B   D   F����   H   J����   L   N   P   R   T   V   X   Z   \   ^   `   b   d   f   h   j   l   n   p   r   t��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       u   ?D�=y�#?%`BD�� D�  >B�\>�jB�  @�     D�� B  BM�>���B�     B�        @��>ě�>gl�>cS�B��=P�`=��#B@  ?.��A�  >�S�B�     D�� ?}�-?�y�L��>���   B���?N��   D�  >�I�@@  @@  @�  >���@�  >%D�� B�ff>�ĜD��       ?3t�>|�D�� B�  >D��@�\�B�b$Bn[q�ʳ�B%{�;�������h>ޑ�A��dBa.��A��C�r���;B~aW��U9BFTt�,�PB��ߟB�MA�@*� #H@�DB~����N]A��2DAv�Bu��z'�A��7��l A>ۧBN	�A0k4B�*�¶2���}VA_���Z��B_B�+PA���;�!û9��������6�4��A���B��C���qo?�M�L       split_indices[$l#L       u         	            	                                                           	   
                                             	          	                           
                 	         	                                                                                                                                                                                                                                L       
split_type[$U#L       u                                                                                                           L       sum_hessian[$d#L       uE�8 EC0 Ew@ E7� C4  B�  Eo� E� D	� A�  C  B`  Bt  D�� E/ D�  C�� C�� BD  A0  Ap  B�  BH  BP  @�  A   BT  D @ D@ D�� D�� D�` C  C  C�  C�  ?�  A�  B   @�  @�  @�  A  A�  B�  @�  B,  B  A�  @�  @@  @   BL  C�  B�  C�� A�  D4  D;  AP  D�  D�  A0  A�  B�  B�  B�  C*  C  C�� B�  @�  A@  A�  AP  @@  @�  @@  @@  ?�  A   @@  A�  BL  B  @�  @   B  A   A�  Ap  AP  @@  @@  @   ?�  @   ?�  ?�  A�  A�  Cd  C8  A�  B�  C�  CW  ?�  A�  C  D� C�  C�  A@  ?�  AP  D�` L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       117L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       G>8S2>���-��F�A$)������`Q�������BtU��^z�hIB4��NU@�����6A S�C#��G�B�������?�U��fLXB�|@3��C�N�C$�CÉ��B!���d#�C�@BA�C��?�5���C$�qB�U�?p��A��7�'�!B>^"���@@����5ْC&O�T���yZB��� ^��%A�u��A���c�����B|M�C}j��z��B)G:�C]B	��h��¿sr��&��$?B�$�A���B���@�@�Q��yL       
categories[$l#L             	                            	   L       categories_nodes[$l#L                      "L       categories_segments[$L#L                                    	       
L       categories_sizes[$L#L                                          L       default_left[$U#L       G                                                                 L       idi;L       left_children[$l#L       G            ����   	   ����                  ����               !����   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E��������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       GG���H�T�H gHHz�    I-��H�0�    H�>IR��I��tI
`1H��G���    H���I�BI���J��H��"    I��H�ՖG��;H�H�XI��H��XI�MqI*�H��I��I���GL~�H�X I0��Hu!�IH~H���                                                                                                                                L       parents[$l#L       G���                                               	   	   
   
                                                                                                                             !   !   "   "   #   #   $   $   %   %   &   &L       right_children[$l#L       G            ����   
   ����                  ����                "����   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F��������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       G>8Q�>�+>;dZ@@  �F�B�  >?|���`Q   B|  >��>�I�=�FBF  NU@�     >hs>B�\=��-B���D�� =��#B  B�33@�G�   D�  >�=q?G�>�t�   >u@�     >x��>�$�>�=q?�(�A��7�'�!B>^"���@@����5ْC&O�T���yZB��� ^��%A�u��A���c�����B|M�C}j��z��B)G:�C]B	��h��¿sr��&��$?B�$�A���B���@�@�Q��yL       split_indices[$l#L       G      	                                    	                                 	                                                                                                                                                                                  L       
split_type[$U#L       G                                                                  L       sum_hessian[$d#L       GE�8 A�  E�` A�  ?�  D�� E�� ?�  A�  Df� C]  B   E�� A�  @�  D]� B  C  B�  A�  @   D1  E�� @�  A`  D\� @@  A   A�  C  A�  A�  BH  A   A�  D&� B(  B  E�` @@  @�  A   @�  D*  CK  @   ?�  @   A   A�  A  B�  Bl  @�  A  A�  @�  Ap  B  @�  @@  A0  A0  B�  D  A�  A�  A   A�  D7� E�p L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       71L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       o=���G�?�;������A� ��:��*�cAhCҋ�?�AW�C.���
��'����B��B:s�7J�B��SA����=��C���RBq�`C����X���B�BDB��������iB�k�C�����@BT�T��x/��e,B:q�Bn?�����d��ûq�C����1[C,�����;CC��A}W�A��C�	B����pA�����.��CUåpVC3�H�J�!�������B>���DB>����@��gC�j@�Y�¬�B;�A44��t�B�~�A��4�2�3B4 ���@A��@u�4¡D�@��"�-�u�o]C�-@�4���A̯��"$�B�w5BYV��1ԗ@/B���A�/�������BB��pC'���Ba'?��n�Q��.����8B�RN?��gA@����?��B���L       
categories[$l#L       -                    	                                     	   
                           
                               	   
                    L       categories_nodes[$l#L       
                        /   0   8L       categories_segments[$L#L       
                                                         *       +       ,L       categories_sizes[$L#L       
                                                                      L       default_left[$U#L       o                                                                                                     L       idi<L       left_children[$l#L       o               	                                    !   #   %����   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M����   O   Q   S   U   W   Y   [   ]   _   a����   c   e   g   i   k   m��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       oHAI@xDH��7H�N�I,�{I�6�H�]�II�G�w�IT�TI6%6IG�<H܁IE��I_�$IRc�H��I J    F���I�
�H��OI*�I��xI�8H���I?��Iz��Hh�8HF(I		�I��H|�pHԪhH脬H��<I8�;I��E��R    I��I�O�H M�G?��Hf��H�:I�U�I��G��yH��    H ��H�s�IyI;��HKC`G���                                                                                                                                                                                                                    L       parents[$l#L       o���                                                           	   	   
   
                                                                                                                                   !   !   "   "   #   #   $   $   %   %   &   &   '   '   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   4   4   5   5   6   6   7   7   8   8   9   9L       right_children[$l#L       o               
                                     "   $   &����   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N����   P   R   T   V   X   Z   \   ^   `   b����   d   f   h   j   l   n��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       o?}p�@�  ?���      B�  B�  >   ?L��=�S�?��>�9XD�  B�  >�dZ?aG�      >s�FB��S      ??}   >׍P>�Q�>XbBp  ?�?�(�> ĜD�  >�jB33?E`BB<  >�@�  >��@�  ���>t�@�  Bճ3>�=q>R�=�v�      >{�m?�{B���B�  Bf  =�t�=Y�   A�  �J�!�������B>���DB>����@��gC�j@�Y�¬�B;�A44��t�B�~�A��4�2�3B4 ���@A��@u�4¡D�@��"�-�u�o]C�-@�4���A̯��"$�B�w5BYV��1ԗ@/B���A�/�������BB��pC'���Ba'?��n�Q��.����8B�RN?��gA@����?��B���L       split_indices[$l#L       o                                                            	                                 
      	            
            
          
         
   
            
                                                                                                                                                                                                                                              L       
split_type[$U#L       o                                                                                                     L       sum_hessian[$d#L       oE�8 DG� E�@ D5@ B�  D� E�0 CU  D   A   B�  C�  B8  E�� A`  C  Bp  C�� C  @�  @�  Bd  A  C�� CI  A�  A�  E�h B,  @�  @�  B�  A�  @�  BT  C�  B�  B�  B@  @@  ?�  B  A�  @@  @�  A�  C�  BD  C  @�  A�  ?�  Ap  E�� A�  B  @�  @�  @   @�  @   A  B�  A�  A  @   @�  BD  @�  B  C�  B�  @�  A�  B�  A�  A�  ?�  @   A  A�  A`  A  @   ?�  @�  @   @�  AP  A   C�  A�  A�  B�  B�  @@  @�  A�  @�  A`  ?�  Ev� D�  @�  A�  A�  A�  ?�  @@  @   @@  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       111L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       K>o����W?E!��8���>�?]EB�|zC�5����7��A�0��^u�?�0gB����ƋIA���B�f�|}�r��_��bV���o�B�oc� ��A��Am1l�#��B^�M�4�3Aj�-�'`AHG~H��$eA�e��x[��	�lA��+B%7>�/¼��$ �B_����>B Y�$��V�@��4A�X@AI�������Bg�5����{���V��3AS�?�Lg���?Bz���q��`�������>5C	&�AV���Z#�>b�B3ml@��~�_���N��?"�J�վ�L       
categories[$l#L                            	                                           	   
                  L       categories_nodes[$l#L       	                  #   %   -   .L       categories_segments[$L#L       	                                           	                     L       categories_sizes[$L#L       	                                                               L       default_left[$U#L       K                                                             L       idi=L       left_children[$l#L       K               	                        ����      ��������      !   #����   %   '   )   +   -   /������������   1   3   5����   7����   9����   ;   =   ?   A   C   E   G   I����������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       KH,Hy�pH9_H0HM��G�ɒH���G�0FH ?�G��Gc��I!
�HJ`�    G��DE���        Hq�G, IEX�     FO8I>��I�Z�H�tZH�!�EqP            H8�
H�%E���    C��     B�7P    IE�IZv�H�^IIa�I2@�I��=G��lH�i\                                                                                                                L       parents[$l#L       K���                                                           	   	   
   
                                                                                               !   !   #   #   %   %   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .L       right_children[$l#L       K               
                        ����      ��������       "   $����   &   (   *   ,   .   0������������   2   4   6����   8����   :����   <   >   @   B   D   F   H   J����������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       KA�     A�  @   @�  >��@�  >���=� �>��A�  @B�\>;dZB���      B�f�|}>���   @   ��o�A�     D�` ?7K�<49XBDp��4�3Aj�-�'`>�l�@o�PA�  A�e�   �	�l   B%7@�  @�  ?<�@E�=�%>bN      @��4A�X@AI�������Bg�5����{���V��3AS�?�Lg���?Bz���q��`�������>5C	&�AV���Z#�>b�B3ml@��~�_���N��?"�J�վ�L       split_indices[$l#L       K                   
         
                                                                                                                       	   	                                                                                                                      L       
split_type[$U#L       K                                                                  L       sum_hessian[$d#L       KE�8 C  E�� B�  A�  E�p A   @�  B�  A�  @�  D@ E�� @�  @�  @�  @@  @   B�  @�  A@  @   @�  C�  CS  D�@ E�x @�  @   @@  ?�  B�  B   @   @   A  @@  @   @   CK  C  A�  C;  C� D� Ap  E�  @   @   BX  A�  B  @@  ?�  ?�  ?�  A   ?�  ?�  C-  A�  C  A0  A   A�  @�  C7  A�  C� B�  C� A0  @�  E�( C�� L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       75L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       C=�G�>\����@�=5�k�@I�4������BBj���6�A��Ad��՝>��YB�$��1��UPB�û��<iB�Y@�yì%������c0A��CH�h��§yw����Õ�'��8�B�0M�Z^��S-B�Yÿh"�B�@��=��|�,Au�$��A�]4��@�»�b�lrOA\��C�4A��ϦB�|�A�TF��{@��q��0���hWBw����B8��Bm)@�����ԡ�|�`�<�M?���<.�BQ��L       
categories[$l#L                  L       categories_nodes[$l#L                "L       categories_segments[$L#L                             L       categories_sizes[$L#L                            L       default_left[$U#L       C                                                             L       idi>L       left_children[$l#L       C               	��������                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A��������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       CG�ԋG�4:F� �I5?H���        I v�Iٔ_H��Is I}BI.@I%(I���Hټ�I��Ie�\Iq��I��I>`�Hw�TI8|H�ۖH�+�JMEI���H˚�H���I2�NI� JI��I9þI�
3IԬ                                                                                                                                L       parents[$l#L       C���                                               	   	   
   
                                                                                                                                         !   !   "   "L       right_children[$l#L       C               
��������                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B��������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       CCB  ?
��>��7>��B$  @I�4���   ?�B  D�� =�S�   =o? Ĝ?�=q>��>�7L?�7D�` >ۥ�>T��<�C�B.  BL  ?���>��m=e`B>49XBճ3@�  >�7L>��`?4�j   �h"�B�@��=��|�,Au�$��A�]4��@�»�b�lrOA\��C�4A��ϦB�|�A�TF��{@��q��0���hWBw����B8��Bm)@�����ԡ�|�`�<�M?���<.�BQ��L       split_indices[$l#L       C         
                                      	      
   	                           
                  	                                                                                                                                      L       
split_type[$U#L       C                                                                L       sum_hessian[$d#L       CE�8 E�� A   D�� E� ?�  @�  D�  C�  E�x C�  Du@ D"� C+  C3  E�x C@  Cl  Cf  C  DO  @�  D!@ A`  C  C(  A0  B�  E�h A�  C/  C;  BD  CB  B  B�  B�  D6@ B�  @   @�  B  D  @�  A   B�  B�  A�  C  @�  @�  A0  B\  D  Ep� A`  @@  C  B  B�  B�  @�  B4  B�  C   @�  A�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       67L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       s���s�/��@ȩ�>����^�A�?R���4��\]B[
c��th�><\@��Bg^���qA�Lj@髭�[�B$��C2n_A�+��Z5�òحYq�B�B��Cz�A�����JA�s4��N�@&S�B����d�?�y���?=B���B0�j�5pW��pbBq����-BX.�.�C-(@ˇ9­m�C����RBԼ�C�7��B�S���?zB;��¬���>L�BOwA��οOh���7Bm{@Y������Be�"����B�[���v��A���A��������@��4@�"|�Ry��a{B��Aj���*����d�BO�W�Y�� �aC!�@�g�9(�B,�CA`eM�`�wBq;�����A�M·�tBAF��C;MJ��J¸���XA���C7)��[(�B�a-��F�@�Z�r��B�x�-��c�����2BK�AFpBv��L       
categories[$l#L       #                                    
         	                         	                               	   
         L       categories_nodes[$l#L       
                	          *   /   2L       categories_segments[$L#L       
                                                                       L       categories_sizes[$L#L       
                                                                      L       default_left[$U#L       s                                                                                                  L       idi?L       left_children[$l#L       s               	                                    !   #����   %   '   )   +   -   /   1   3   5   7   9����   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c   e   g   i   k   m   o   q��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       sG��I;�ID�H���I�3�IKR�H���H��I�� I�Iv�\I� IץRH�wzH�-�I8��I��^H���    I*rI���IYBpI��I�/I�?I�Iq	�IV�H���H�N�    I/w�I�YpIj�~IE�H�H�HƸ�H�B�G�]|IA <I�RIrh�G���IY�H��IZ�Iw��H��HF��H��@I�b�IV�I���IbQ�H��UIΖH�e4H�͏H���                                                                                                                                                                                                                                L       parents[$l#L       s���                                                           	   	   
   
                                                                                                                             !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   :   :L       right_children[$l#L       s               
                                     "   $����   &   (   *   ,   .   0   2   4   6   8   :����   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d   f   h   j   l   n   p   r��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       s         ?L�D   >���@@  >�7L@�     @�  ?%�>��`?��!A   >��7>\)B.  C2n_@�p�?�-@d��@L(�?4��A�  @�     =#�
>�Q�@�  ��N�D�     =Y�@   ?N�?!%?���>�!?��@~{>��w   B@�@   ?!��B.     =� �?K�   >��PB�  Bj��>�v�?��>�\)?��?�PA��οOh���7Bm{@Y������Be�"����B�[���v��A���A��������@��4@�"|�Ry��a{B��Aj���*����d�BO�W�Y�� �aC!�@�g�9(�B,�CA`eM�`�wBq;�����A�M·�tBAF��C;MJ��J¸���XA���C7)��[(�B�a-��F�@�Z�r��B�x�-��c�����2BK�AFpBv��L       split_indices[$l#L       s                                       	                                                    
                            
            
                                            	      	                                                                                                                                                                                                                                   L       
split_type[$U#L       s                                                                                                         L       sum_hessian[$d#L       sE�8 E�  Ep E�h Cɀ D�  D+� E�@ C%  C�  BD  D�  C�  C�  CU  E� D�  C"  @@  C*  C8  A�  A�  D|  B@  C  C�  C�� C?  CR  @@  E� C*  C�� D�� Bt  B�  C  A`  B�  B�  A�  @�  A�  @�  Di� B�  B(  @�  B�  A�  C2  B�  B(  Cq  A�  C+  Bh  C  CB  E� B  C  C  C�� A�  D�@ AP  B@  A   B�  C   A�  A@  @   A�  B�  B  B   @@  AP  @   @   A�  @�  @   @�  D^� B0  B   B(  B  @�  @@  @@  B�  @�  A@  @�  A   C(  B�  @�  B  @�  Bt  C4  Ap  @�  B�  B�  BT  @�  C  A�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       115L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       i=�E?Y����?�ޠ���T��A���?���B�_���>A�B�C\<�v&�Cb*�A4g$>~�B-C*��C ���B��{B����PC�~�@�'�����TS�W�C�7��k��Bn?4�,��jB�rx���]A�,�C�^��( Á��V��?5CC���D��|�CW�k�.O B6B�B�|-A�Z�BDB;�|B��S�B-'��oӳC
�A��TCa�»��C,�����>����܊?���5H�B��YA�?���eµ��A��K�9�lC3FA��~r�AzzM���!º}z���6g@����\��An�gBJ���UP`A���A��B�YzAW ���'�1A��9�O��B�L���AƆQ�_�³�8B�S7@ϏgA�k��&B�	MAA#QB=C�K�\L       
categories[$l#L       -                                	   
                              	             	                                            	   
                  L       categories_nodes[$l#L                                        %   '   ;L       categories_segments[$L#L                                                                                     *       +       ,L       categories_sizes[$L#L                                                                                                  L       default_left[$U#L       i                                                                                           L       idi@L       left_children[$l#L       i               	                                    !   #   %   '   )   +   -   /����   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q����   S   U   W������������   Y   [   ]   _����������������   a   c   e   g��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       iG��H�y\H�m�Hd�NH�amH�jH� �H��
I*�Hp��HzD<G��H�-�H��tH�q�H��]I�oI���Gġ0H�G�@2H �H>�GtJ�    H�dMH�IpH,��G�8HڂtI3t�HE|SHF.rIP�H���H�0I�F,�2Fa� G��8H�E�@�    F`��E��Gm            H���H��lH��HK�                G�TH��3H�X�H�U[                                                                                                                                                                                L       parents[$l#L       i���                                                           	   	   
   
                                                                                                                                   !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   +   +   ,   ,   -   -   1   1   2   2   3   3   4   4   9   9   :   :   ;   ;   <   <L       right_children[$l#L       i               
                                     "   $   &   (   *   ,   .   0����   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R����   T   V   X������������   Z   \   ^   `����������������   b   d   f   h��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       i?pbN?��@D�?}�      @H��?KC�?N��@��HBH��      B8Q�@@  ?���@X           @@  >���?��R@�  @�'?�ȴ         D�@ @�  ?q�B8Q�@@  @�  D�` @�     D�     D�� BD  ��D@�  B  >�33B6B�B�|-A�Z@�  B8Q�?e�B4(�B-'��oӳC
�A��T@@  B
ff   D�� >����܊?���5H�B��YA�?���eµ��A��K�9�lC3FA��~r�AzzM���!º}z���6g@����\��An�gBJ���UP`A���A��B�YzAW ���'�1A��9�O��B�L���AƆQ�_�³�8B�S7@ϏgA�k��&B�	MAA#QB=C�K�\L       split_indices[$l#L       i   	                     	   	                                          	             
                                                                                                                                                                                                                                                                                                   L       
split_type[$U#L       i                                                                                            L       sum_hessian[$d#L       iE�8 E�� C�  E�H BP  CA  C)  E�� B(  B  A�  @�  C<  A   C!  E�h C  B  @�  A�  @�  A0  @�  @�  ?�  B�  B�  @�  @�  B(  B�  E�H B  B�  B  A�  A  @   @�  A�  A@  @�  ?�  @�  @�  @�  ?�  @   @   A�  B(  B�  A�  @   @   @@  ?�  @�  B  B  B�  E�� A�  AP  A�  Ap  B�  A�  @�  A   A�  @�  @@  ?�  ?�  @   @@  Ap  @   @�  @�  @   @   @�  ?�  ?�  @�  ?�  @�  A�  A   A�  A�  B�  Ap  AP  AP  @@  ?�  @�  A�  A�  A�  A0  B�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       105L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       A=��>N�η?ƤF�1Tv?ۻB�
y��,�Bp�R?�AQ��<X�&S$Cc}.A����'�VC0W��6>��B�[ÕC#;� ?^C�C��D��B��[��p����� �B���C�VA�xÙ�S?��u��A���1�����������gC �@�i���9@F\gCL�3�LqB{��B�AC~��ByNL@�h�B�i����
/AM�N#����B@��g��B)� C5<��Hb�A����'W����L       
categories[$l#L             L       categories_nodes[$l#L          L       categories_segments[$L#L               L       categories_sizes[$L#L              L       default_left[$U#L       A                                                          L       idiAL       left_children[$l#L       A      ����         	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?��������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       AG�~gGژ�    H��0I�4H�I��#InI1ZHE�J<�I��*I���I���I}R!IN�IlH�o�I��I��XI�S�I�O�I���I'�I
g�I��BI��PIivI�ƾIPHIF��C\�                                                                                                                                 L       parents[$l#L       A���                                                     	   	   
   
                                                                                                                                      L       right_children[$l#L       A      ����         
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @��������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       AA�  B�  ηB�  D�� B�  D�  >�o?>5?B�  >��>�o@�  >1&�D�  >��A
=B�33>��@�  A�  >o@�  >q��A�  A�     >��\>��>���?�=q?�-B̊=?��u��A���1�����������gC �@�i���9@F\gCL�3�LqB{��B�AC~��ByNL@�h�B�i����
/AM�N#����B@��g��B)� C5<��Hb�A����'W����L       split_indices[$l#L       A                                                                                      	                                                                                                                                               L       
split_type[$U#L       A                                                                L       sum_hessian[$d#L       AE�8 E�0 ?�  EĐ DE  E�� B�  D,@ B�  E�p B4  BP  B  CV  C� B  B�  E�0 C  A�  A�  A�  A�  A�  @�  C$  BH  C�� B�  A�  A   Bp  @�  E�  C"  B�  A�  A   Ap  Ap  @�  A�  A`  A�  @@  @�  A�  @   @@  B(  B�  A�  B   C  CR  @�  B�  A�  @�  @�  @�  Ap  B4  @�  ?�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       65L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       {=��N���@�A&D���bھ�&
B��7x�A��r�B���G��?�U�§0A�v�C��pAd�¦/B��QA@[ �����U���
xB.��B��BĀ`��f1C0�A�̣�''B��DR}�A��W�A!"B���̦�n��C
��C`_.@�i��uB���B��?�KCAe�Kh%CI���?2���#�A��D
)�C5}�#�#Cw�7�3A�9.C����=�ïʦCkv��Z�B�B�C���@}��C�4B�+�������~�B�Y*��[�����A��;�ĿB��cA�;D�.��B������K@��´��A����h²�tC]�)�����)A�G�AF�y��>��ιNBm�B�i@t�aB��i�O�?,�v�x���(s�Cd�B.����5�C�,�B*�@���C ��S��B�6@��B�'���AM4��Q�AH��C6��A���A��s�����G�B�MRA&"��'B��L       
categories[$l#L       :                                         	                                     	   
                                             	   
                                     	   
             L       categories_nodes[$l#L                         !   #   $   )   6   8L       categories_segments[$L#L                                                                "       +       8       9L       categories_sizes[$L#L                            	                                   	                     L       default_left[$U#L       {                                                                                                         L       idiBL       left_children[$l#L       {               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c   e   g   i   k   m   o   q   s   u   w   y��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       {G��H��HҥjH���H�m�I��I�bI
��I�$I.r�H�mmI I�I@vI,��J�dI1h�I��IP�H�FuI���H���I��I\�~H��I�
�Izh�H�űI���I1��H�+I_I��I��I8I�~H:��H�-�Hw�H��sI3�<H�L/I���H���H�ɶH�_�I�n:I" H�tI��I=)�IK{H�H��<G�&8F�]�IEfI3'H�/*H}��G�g�HXU�                                                                                                                                                                                                                                                        L       parents[$l#L       {���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <L       right_children[$l#L       {               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d   f   h   j   l   n   p   r   t   v   x   z��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       {A  D�� >޸R?   >�hs>�?K�>�\)??}?@  @Ĝ>��;?M�?ǍPB[��Bճ3      >š�D�� ?o\)      >�ƨ@�H   A   ?f$�B~?)�^A@  B̊=>A�7   @>{      >��7?���>� �?*=q   A (�@�  A  >\>�A�A��?@  D�� D�� >ڟ�D�  B'
=   >�\)   ?Z@   ?�^5@�G�B�B�C���@}��C�4B�+�������~�B�Y*��[�����A��;�ĿB��cA�;D�.��B������K@��´��A����h²�tC]�)�����)A�G�AF�y��>��ιNBm�B�i@t�aB��i�O�?,�v�x���(s�Cd�B.����5�C�,�B*�@���C ��S��B�6@��B�'���AM4��Q�AH��C6��A���A��s�����G�B�MRA&"��'B��L       split_indices[$l#L       {            	         	   	   	   
         	   
                
      
                             	                                   
                                              
                                                                                                                                                                                                                                                                       L       
split_type[$U#L       {                                                                                                                L       sum_hessian[$d#L       {E�8 DՀ E�� DX� DR� E�� CÀ C�  C�  C�  C�  E�� B�  C�� A�  C�  B�  B�  C�� B�  C�  C�  C*  E�0 BX  B�  A@  C�� A�  A�  @�  C�  A�  A�  B�  A�  B�  A  C�  B   B�  B8  CV  C-  C  Bt  B�  E�0 B   B@  @�  A  B�  A   @�  C�� A   A�  A  A0  @�  @   @@  C�� ?�  @@  AP  AP  A   A@  BT  @�  A@  A�  B8  ?�  A   B�  C�  B  @�  B�  @�  @�  B  C:  A�  C	  B  B�  @�  A�  B  @�  B�  E�� C	  A�  ?�  A�  A�  @@  @@  @�  @@  B�  ?�  @   @�  @@  ?�  B�  C�� @�  @�  A`  @�  @�  @�  A  @   @�  @   L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       123L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       5>�}'?!o��)>�>;C�@���4���?�O��Cba�*�������%�?V�������B}z�B�P�u�4@d���C>B�A���ç��?5[�C��A��g°�A�m@�$g����?�镾��3C�m�����B����C��4��v8>��B�j@�JA�	����4�z��tA˪��y�AA���f�C@�A��L       
categories[$l#L                                       	   
                                            	   
                    L       categories_nodes[$l#L          
               !L       categories_segments[$L#L                                                  L       categories_sizes[$L#L                                                 L       default_left[$U#L       5                                                L       idiCL       left_children[$l#L       5               	   ����               ����         ����   ������������      !   #   %   '   )����   +��������   -   /   1   3������������������������������������������������������������������������L       loss_changes[$d#L       5G��^Hw�H��"H2��H�*fH��`    H
2�H;�G�TG'�NH��	    I ��HoTG3h    A/l             H)*�H���I	XiHRHG�i;G�	�    E�L�        H<��HM�F��lF~3�                                                                        L       parents[$l#L       5���                                                     	   	   
   
                                                                                         !   !   "   "L       right_children[$l#L       5               
   ����               ����         ����   ������������       "   $   &   (   *����   ,��������   .   0   2   4������������������������������������������������������������������������L       split_conditions[$d#L       5C  C   ?��B�  B�  >����D�` >�hs<�   ?!G����D� B�  =\)���   B�P�u�4@d   D�� >�G�=D��<���   A��g   A�m@�$g@@  =��   @�  ����B����C��4��v8>��B�j@�JA�	����4�z��tA˪��y�AA���f�C@�A��L       split_indices[$l#L       5                  	                    
                                                                                                                                                       L       
split_type[$U#L       5                                               L       sum_hessian[$d#L       5E�8 E�  B�  Eڨ A0  B�  @   E�h A   A  @   B�  @   A�  E٠ @�  @   @@  @�  ?�  ?�  Bp  @�  A�  @�  E�x @�  @   @�  @   ?�  AP  B<  @�  @@  Ap  @�  @   @�  C�� EА @   @@  @   @   @�  @�  AP  B  @@  ?�  @   ?�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       53L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       }>!{@k��a}�?9�$B,A]}��/w�@0��Z�AB�B�d���>�Bj�������?�`YB�f�C(��½2mB5~���`BP��CA�A@�}�´<�A���CD$���{
�q�B˱��s#@9"A��IC���C���ƺ��Ý��z	]C3 ,���c×4i��p�B�}>D	W�B����V_AQ��B$.��@B՞�WC�C���@W�I���B����5�A�'[C��	ޟ�
�l?��?�`<�DA�"��ae�ʥ�A��[BC�C3F�A� �C*v/�̃n�"���������@@ao�£��Av�#B�b-��{B.m������5����{�B��A��B��YB�w�CaOL�V"wBV���y$���t�$��@�!�C*�8��;���DkAS�N��AuL���q��̀|C�>��4����A�v��F�A?�RC��A��g��%B.�B�b��6�gCt+�A�!�@�#�Aq�W�xU�A�%O��L       
categories[$l#L                                   	              L       categories_nodes[$l#L       	   	            "   '   /   2   :L       categories_segments[$L#L       	                                                  	       
       L       categories_sizes[$L#L       	                                                               L       default_left[$U#L       }                                                                                                                L       idiDL       left_children[$l#L       }               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G����   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c   e   g   i   k   m   o   q   s   u   w   y   {��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       }G��H�v�H��PH�խI0�"IYL�I���H� I$x�I
��H�q�ID��I� mI�4�I$9Hx�~I2)�It\I��H���Ip�IV��If��I8��JJ�I+.I�E2IU}JKIᬷI�{HkF�I8p�H���H0��I��    Ho�HS��H�d�H�Y�H��FIjߞI �I�2NH��I�I&�I�I��I�7>I `LHl� I�o IH��H�t$H�]�I���I�9J `�H�vFIOg�I��                                                                                                                                                                                                                                                        L       parents[$l#L       }���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <   =   =   >   >L       right_children[$l#L       }               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H����   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d   f   h   j   l   n   p   r   t   v   x   z   |��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       }@Vff@FffD�  ?�ȴD�� @�  D�  ?N��=� �   A�  B�  B�  B�
==��D�     B�33      B@�>]/@   @Z�HA`  B�aH@�ff>aG�@���>��>�Z@E�>aG�@      A�  ƺ@7
=B     B~>k�>>v�A   BH��BK��D�     >��?O�   =�\)>��7C  ?�h@�  =�9XB�     @�p�?�?$ZD�` ?�`<�DA�"��ae�ʥ�A��[BC�C3F�A� �C*v/�̃n�"���������@@ao�£��Av�#B�b-��{B.m������5����{�B��A��B��YB�w�CaOL�V"wBV���y$���t�$��@�!�C*�8��;���DkAS�N��AuL���q��̀|C�>��4����A�v��F�A?�RC��A��g��%B.�B�b��6�gCt+�A�!�@�#�Aq�W�xU�A�%O��L       split_indices[$l#L       }                        	                     	                                                       	                                                            	   
                        
                                                                                                                                                                                                                                                              L       
split_type[$U#L       }                                                                                                                    L       sum_hessian[$d#L       }E�8 Ea� EX� ER0 C|  D�� E� EL B�  B�  C<  D6@ C�  B�  E@ EJ  A�  A   B�  B   B   C   A�  D@ B�  C�  BX  B�  BL  B`  E� EG� B(  A�  @�  A   @   B�  A  A�  A`  A�  AP  B�  B�  @�  A�  A`  D� BX  B(  Cw  A  A�  A�  B   A�  A�  A�  A�  A�  D� DР EF� A�  A�  A�  @   A�  @@  @   @�  @@  BD  A�  @�  @@  A`  @�  A   @�  A@  @�  A   @�  B�  @�  BP  B  @@  @   @�  A�  A  @�  A�  D� @@  BL  A�  A@  AP  Cj  @�  @�  A�  @�  @@  A�  A�  A   @   A�  A�  @�  @�  AP  @�  A�  A0  A�  B�  C�  B�  D�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       125L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       {>'z�AE��zU��,A�tk@̂�����A骖���B|n��ր@�7@C<.2@��O�X����i6B���A��s��@A B��C�(���['Bt��?)�D����|A��k��n}�->��B����#��p�CXB�7R�"��WS7�p�}���C�<C%<�Aɶ�A,@D7)���MPµ�+�t�%B�v%�z?A<�zB��
C��RB��9�{k;A7B��o�#��A��?Aa��¥�)B&J�3�A�[C<6pB%~@¤�?B����Bk���VB6$�nT�¥�:>�K�A$���Fy��E�¼��BP������B�o7�0,�C���B,���$�"B	0@׾M�w B�׊Cr����%B�F��Z���#�.�B@B�B'A�XN>:���п�5�A(N<��9�BP���w�¾ |����A���B�XA�Kg�����ب�Ay'����A�*K�����[=��@�AO�����l����^�L       
categories[$l#L       '                             	   
                                           	             
                                     L       categories_nodes[$l#L                             '   +   ,   6   :L       categories_segments[$L#L                                                                               !       #L       categories_sizes[$L#L                     
              
                                                 L       default_left[$U#L       {                                                                                                           L       idiEL       left_children[$l#L       {               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c   e��������   g   i   k   m   o   q   s   u   w   y������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       {G�q�II��Hh��I�)dIH�IC��H��I� I�;nIH��I�J�IMJ��I-��IJ�I���I2xVI] |IrS�ImɵIfZ@Im�rH��&IO��H�!�I�m�H֘Iq-*H�I�I�I�AI�6I�9DI	I�*H�1RH��2I�	I2PIC��I}�hI��I��D6pPF�# IF/�H��H鼗Ii�IYz$I�0        HC�~G!��IP�I�@�H�ڔH�äI;�]Iȍ�Ip�H�'                                                                                                                                                                                                                                                L       parents[$l#L       {���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <   =   =   >   >L       right_children[$l#L       {               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d   f��������   h   j   l   n   p   r   t   v   x   z������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       {   >["�>ٙ�>ix�   >׍P@,��>�+   D�  =y�#=��>$�/   ?��>`A�>x��A�     >���@�G�>`A�@�H=,1>Y�@�  D�� ?��>���   >��>^5?>t�?jA  ?Y�#>1'BM�D�     @�@@  @�        ?�I�@/
=>��j=�+>dZD�� B��
C��RD��    ?���=�S�>B�\   @Vff@1G�A��>O�A�[C<6pB%~@¤�?B����Bk���VB6$�nT�¥�:>�K�A$���Fy��E�¼��BP������B�o7�0,�C���B,���$�"B	0@׾M�w B�׊Cr����%B�F��Z���#�.�B@B�B'A�XN>:���п�5�A(N<��9�BP���w�¾ |����A���B�XA�Kg�����ب�Ay'����A�*K�����[=��@�AO�����l����^�L       split_indices[$l#L       {         
          
      
                	          	   	               	                            	   	   
   
                                          	   	                                                                                                                                                                                                                                                                                              L       
split_type[$U#L       {                                                                                                                L       sum_hessian[$d#L       {E�8 D�� E�� C�� D(@ E� EdP CS  C"  C�  C�� EP A�  D�  E� B�  B�  B<  B�  C  CE  @�  C�  C  E	� @�  A�  D0  D@ DR@ D�` BD  B0  Bp  Bh  A�  A�  BT  Bx  B�  B  B�  B�  @@  @�  Cy  B|  B$  B�  Da� D�� @�  @   A0  @�  D� C	  C�  CE  C�� C�  C�  D�  B@  ?�  AP  A�  A�  B  BH  A   A�  @   A  @�  A�  A�  A�  B(  Ap  B�  A�  A�  @   B�  BX  A�  ?�  @   ?�  @@  Cu  @�  A�  B  A�  A   A0  B�  D2@ C>  D8  D  @�  @�  @   @@  C�  C'  A�  B�  C�� B�  C  BT  B�  C�  A  C�� C�  A�  C+  Dq� L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       123L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       o>���@n���F?�S Cy�A�@��p᜿,UB2<C���B�]��>��B�w�O� �/�!�wX@9T���=Bkz?Cm�d������,4c@��<B�La�O��B^������,@�p��e�m�O��AG�IB�/: �C;;�A�98����C���A ����I�hC@b�â��B�Q�A�s�� A�ذC.��=۴��5����jC	ǁ�x��P(B�Aq�7����A�1����5PP������A �ܿ�]�B����@%�"�4�fB�3�A-�pA�T �a�A��a���B!<�B��AJ���ZL�@�Yc��-�B���@�#��(DD��mw���gB.�AԂ���gA\$���Bw,��7��ǜ�B���?�p��E�&�t���A����nC(�`BC�^J�A�f��	}��-
0���B���	�RgL       
categories[$l#L       	                             L       categories_nodes[$l#L                   %   -L       categories_segments[$L#L                                           L       categories_sizes[$L#L                                          L       default_left[$U#L       o                                                                                                     L       idiFL       left_children[$l#L       o               	            ����                        !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M����   O   Q   S   U   W   Y   [   ]   _   a   c   e   g   i   k   m������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       oGɈ�I&�H��LH��I��fI&4HՄ�H�H�I̀    IF�H��}I��H��I[G�IB��I
QIfIl�BH�)(H�V�H�vI/n\H�DwI/��H���I���I�*�I%��H�I��I0۰I`7�Hr,II] I~�G.G� G��    H?�FG��PG��G;i�H�r�H{��IDE�I!$H���I%D
H�ʪI�I��I0	HH�$�IH%0                                                                                                                                                                                                                        L       parents[$l#L       o���                                                           
   
                                                                                                                                         !   !   "   "   #   #   $   $   %   %   &   &   '   '   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8L       right_children[$l#L       o               
            ����                         "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N����   P   R   T   V   X   Z   \   ^   `   b   d   f   h   j   l   n������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       o>�&�>��@   @�>x��>fffB\33@   >�ƨC���>z�HBu�R@�  BH  >ě�>�?}>'�B'
=>�-   ?-VB\33D�` @8�9D�� D�� @�     >�@�     ?+�>޸R>uD�` >���@�   D�� B�aH���@�  =>�  >j~�   D�  ?U�>�  @@  A   >ܬ?���@Z�H>� �>z�HA@  ���A�1����5PP������A �ܿ�]�B����@%�"�4�fB�3�A-�pA�T �a�A��a���B!<�B��AJ���ZL�@�Yc��-�B���@�#��(DD��mw���gB.�AԂ���gA\$���Bw,��7��ǜ�B���?�p��E�&�t���A����nC(�`BC�^J�A�f��	}��-
0���B���	�RgL       split_indices[$l#L       o               
            	                      	         	                                           
   	                                            
   
                  
   	                                                                                                                                                                                                                           L       
split_type[$U#L       o                                                                                                          L       sum_hessian[$d#L       oE�8 E�  D�` E�P A�  C�  D�  E�� C�  ?�  A�  B�  C�� Dc� C�� Dq� Ez� B�  C�  A@  AP  B�  A�  CH  B�  D6� C3  Bl  C�  D$� C�  D�� E` B  B�  B<  CS  @�  A   A0  @   B�  A  A   @�  C  B4  B�  Bd  D@ CR  B�  B�  B0  Ap  B|  Cy  D� B`  CV  B�  D�� B�  D�� D�� A�  @�  B(  B   A�  A�  C  B�  ?�  @@  @   @�  A   ?�  A�  B0  @�  @@  @�  @�  @   @�  BT  B�  AP  B   B  B   A   BD  C�� A�  C  Bt  B   B�  @   B�  A�  A�  @�  A  A�  B  Cf  A�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       111L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       u>`�@�S��]��B�&t@Ww�Ao"���B�_����BWFw?����_�AoP����}A&'���/C# [�S�B��`B��U�k�:�hA��B����.A����a�I�?	�C|#@�osB����!%�Y&CCu���f·�}@�BE|A��rC(�t¦�(@����{����8�Cq��@ڕ���;�B��a�0�A'�B�E� ��A+_��*rc��l�����u7sB� D2�)C��?v�oA��$ޝ�4�g�BuAv2�����A}'����Bj�%BŅ�A�?���Q�A��:�lA+� ���P�B!]�Cv�A��@A��=?�gv��p����B,���nt��J��д�Bv���~A���D���ܝ@�LpAW�\���}B��k�y�����BD<HB"��+�Z�ϼ ¿��Bw���0lC 3�E��C��B0�'A�:iCj	n@-�X���L       
categories[$l#L       %                                     	               	   
                                            	   
            L       categories_nodes[$l#L              	             !   "   /L       categories_segments[$L#L                             	                                   $L       categories_sizes[$L#L                                                               L       default_left[$U#L       u                                                                                                        L       idiGL       left_children[$l#L       u               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =����   ?   A   C   E������������   G   I����   K   M   O   Q   S   U   W   Y   [   ]   _   a   c   e   g   i   k   m   o   q   s������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       uG�H��H,¦I ��H�Y�HѕaI��H�&�H�RH���H��DIN��HթaI��jI��H�?�IqTH)ްE��XH��4H�I�LIH2H.@�H�N�I3�I���I/7=I�(I�v�II�    G�΀F���I:=ZF��            Hy
�H��p    H6�IlIW TI#� H㈢E[߀H�ZI2*H���Ib��H��zI9�ICz�I ��Ij�2I�XH�IF�I>�I�jIE�z                                                                                                                                                                                                                        L       parents[$l#L       u���                                                           	   	   
   
                                                                                                                                   !   !   "   "   #   #   '   '   (   (   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <   =   =   >   >L       right_children[$l#L       u               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >����   @   B   D   F������������   H   J����   L   N   P   R   T   V   X   Z   \   ^   `   b   d   f   h   j   l   n   p   r   t������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       u   =y�#@�  ?�O�>B�\=���>]/>B�\@j��   >|�   >�\)>:^5>_;dA�  =49X>�(�@@  >׍P@   =�t�>~��D�` >�ƨ   A`  @�>�/>�X=�C�B��         @�=q·�}@�BE|>9X?K�¦�(>���=�\)B\  AP  =o   =�j>�$�A�  @�  >��#@$(�>$�C  >P�`>�I�?�=q>L��D�  B�  B�ffA��$ޝ�4�g�BuAv2�����A}'����Bj�%BŅ�A�?���Q�A��:�lA+� ���P�B!]�Cv�A��@A��=?�gv��p����B,���nt��J��д�Bv���~A���D���ܝ@�LpAW�\���}B��k�y�����BD<HB"��+�Z�ϼ ¿��Bw���0lC 3�E��C��B0�'A�:iCj	n@-�X���L       split_indices[$l#L       u      	                            	                      
      
         	                      	                                       
                                      
            	   	                                                                                                                                                                                                                                       L       
split_type[$U#L       u                                                                                                             L       sum_hessian[$d#L       uE�8 EC0 Ew@ B�  E>� Dv  E9� Bp  A`  B�  E6� B�  D^� D�� D�� A�  B0  A   @�  B�  Bl  D�@ D�@ A�  B�  D� C�� D�  C.  A�  D�` @@  AP  @@  B$  @�  @�  ?�  @@  A�  B  ?�  Bh  CD  D]� A`  D� @@  A�  B4  A�  C�� C~  C�� B0  D�@ B�  B�  Bp  A`  @�  B  D�  @   A0  ?�  @   A�  A�  @@  ?�  A�  @�  A   A�  A�  B  C>  @�  DR@ B4  @�  A  Bt  D�� ?�  @   A�  @   A�  A`  AP  A  C�� A�  B�  C+  CE  B�  @@  B$  DȀ A�  A`  B�  B�  A�  Ap  B4  @@  A0  @   @   B   @   Dn� B�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       117L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       {>{��@
^�b�A��Y�RDZ�YQ������XA��k� �A��A�s�¸�1?���	��I<��uAWf|BuXz�r/A� 0�C�ӕA�D�Cb��@7W7�;a��tq�A��KŨê(AQ[��aIZB���Â���%B.����ԈBv�C�W@s���s�b���0@]( CW�A<s�C��C|2Bs��x��Cu�xB9m(+E��ô�vA���C��<B_ ��C��U�A�D�2�B�����f�A����p�Aֲ���$k��� A�<�r=@���Bi���n�@˭�?��vB� �J�gBk���V�@���L[���&cA�}j����V>���AH������A%1���C�pA6D&@]%�A�6�Ah;���B�zAT�4A酅��	A9Gx��o�B� ��I�!�~J�@�'�B�"��B9�C��JAo_��O#�� �������GZ�F�1��jBS��@�� ��B�<.�"?nL       
categories[$l#L       =                      
                                               	   
                                                   	   
                                                
                  L       categories_nodes[$l#L                            +   .   0   1   2   ;   =L       categories_segments[$L#L                      
                                                 +       ,       -       :       ;L       categories_sizes[$L#L              
                                                                                    L       default_left[$U#L       {                                                                                                   L       idiHL       left_children[$l#L       {               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W����   Y   [����   ]   _   a   c   e   g   i   k   m   o   q   s   u   w   y������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       {H Q@H|O�H�(H�dHhP�H��H��H��dH���H�?jI�xH_�<ID�,H�[�I@�fH��#H�)�H��:H���H�:8I<�4IT\�H��HfiHxN�H��I4��If��H��I[�H�W�Hv��H#}H
��G�}H��lH�c�H�H�-DH�B<I$2If�+I+�DF2pD    H��HQ�    E�1�He\F�0H,��HLFH�|?H.n�I��I�]�H�QpH��`H#8G�7�G�^�H��                                                                                                                                                                                                                                                L       parents[$l#L       {���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   -   -   .   .   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <   =   =   >   >L       right_children[$l#L       {               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X����   Z   \����   ^   `   b   d   f   h   j   l   n   p   r   t   v   x   z������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       {>��   >��@�?d�/>A�7Bճ3>��y>���?+�?f$�=o      >� �   D�  >� �@�  ?�y>�&�   Ap  B�\>�l�@   B4(�B�=q   @�  B�  >���=�/?�oAp  >�\)D�  A@  >�+>���>�bN@�  @�G�   CW�B�     C|2         ?LI�?�  >���D�� @�  @@  D�  @�     B�     D�  ��f�A����p�Aֲ���$k��� A�<�r=@���Bi���n�@˭�?��vB� �J�gBk���V�@���L[���&cA�}j����V>���AH������A%1���C�pA6D&@]%�A�6�Ah;���B�zAT�4A酅��	A9Gx��o�B� ��I�!�~J�@�'�B�"��B9�C��JAo_��O#�� �������GZ�F�1��jBS��@�� ��B�<.�"?nL       split_indices[$l#L       {          
                                                                    
                           
                                                                                                                                                                                                                                                                                                                                              L       
split_type[$U#L       {                                                                                                              L       sum_hessian[$d#L       {E�8 E�� D�� Dy� E�� C0  Dw  C�  D  E�� Ce  Bl  B�  Dp� A�  C�  A�  C�  Cp  E�� C�  @�  C_  @�  B\  B�  A�  C�� D@ A  A�  C�� BD  A   A@  CQ  C7  CC  B4  E}� C�� C�  B(  @@  @@  C[  @�  ?�  @@  BP  @@  A�  B�  A  A�  C�  @�  B�  D� @�  @�  @�  A0  C�  A�  @@  B8  @�  @   @�  @�  C)  B   B�  B�  C  Bp  A  B  E(� D�` A�  C~  B�  C4  B   A   @   ?�  C/  B0  @   @   @   ?�  A�  A�  @   ?�  A�  @�  A@  B`  @@  @�  @�  A@  C�� @�  @�  @   B�  @�  C�  B�  ?�  @�  @@  ?�  @   @�  @�  @�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       123L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       {>`���|?��2A��}�� +B��?Q��?�m�B�\8�0��]�B����)�n�<�W?���­�[A�1C�t�{���B����K%=��.��"�B�IyB}��}�C�V@�$��>0B@�WJ�Ω�ã�!B�[z�A�DoB|ܘ@�@��˪���A�C���A�l���z.B����JpØ��Bo��ÖO�Cs��B��RB�7RD@�u����e��6��-Ia]C�l@2̓�A��e�K@�(�A�ZA�������@�x�B��`��5tAa�CcqBp���αB~����B����B®v���ɵB\�OC<�l��z���B%���3��?��wB�As�u A�a��lmG���B:���$AAdQ�B��A���>���BX�'��`Bg��@Xś�(К¤�=̎��Ь± J�ÑX�vL
BH�?�߭�9@K��ϟB�-i�%}+A��4?Ai�AW����X�Ⱦ�>�S^L       
categories[$l#L                                 	                                       	    L       categories_nodes[$l#L       	                     -   4   7L       categories_segments[$L#L       	                      	       
                                   L       categories_sizes[$L#L       	                                                               L       default_left[$U#L       {                                                                                                            L       idiIL       left_children[$l#L       {               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K����   M   O   Q   S   U   W   Y����   [   ]   _   a   c   e   g   i   k   m   o   q   s   u   w   y������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       {G�k�H�)�HZ�VH���H��I@�6HnMlH��I�H�
�Ij_�Ic8�H6?IM�cH?�&H�Z�H�ВIc�H�c�H�e I�CIM\XIUO0I�PI�XHt�H \I'ӢIW�I-�:H嚄H�H�HXTI��H�3@IZOH&��H��u    I��I5I7��H�lH��TI=�G�H�    G�NuH�$I�^I�G���F�gH+�H6�I
\�HH��xI-�I,wQIt �I@ٴI1E                                                                                                                                                                                                                                                L       parents[$l#L       {���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   $   $   %   %   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <   =   =   >   >L       right_children[$l#L       {               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L����   N   P   R   T   V   X   Z����   \   ^   `   b   d   f   h   j   l   n   p   r   t   v   x   z������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       {>$�D�` >n�   =��#   >�u>2-   =�F?�o>\)>��H>��+=�;d>&�y>	7L?r�>��>��!=���@@     >hs>hsB��{      BV  =�v�=�^5>-V@@  =��>cS�D�@ @�  >D����˪>���@�  @�  >�=q>T��>aG�   Ø��B<=q>��F>�I�>�/Bb     <e`B>y�#   >���?r�!@@  >��\>��H?WK�=ȴ9�(�A�ZA�������@�x�B��`��5tAa�CcqBp���αB~����B����B®v���ɵB\�OC<�l��z���B%���3��?��wB�As�u A�a��lmG���B:���$AAdQ�B��A���>���BX�'��`Bg��@Xś�(К¤�=̎��Ь± J�ÑX�vL
BH�?�߭�9@K��ϟB�-i�%}+A��4?Ai�AW����X�Ⱦ�>�S^L       split_indices[$l#L       {   	      	      	       	         	   
   
      
            
                                                  	                            
                                                      	   	                                                                                                                                                                                                                                                      L       
split_type[$U#L       {                                                                                                                  L       sum_hessian[$d#L       {E�8 D�@ E�� Cy  DN@ CC  E�� CK  B8  D3  B�  B�  B�  B�  E�X B  C)  A�  A�  D*@ B  B�  @�  Ap  B�  AP  B�  A�  B�  D`@ E�P A�  @�  BH  B�  A   @�  A�  @   D  C  @�  A�  B�  A�  @@  ?�  @�  A   A�  B�  A  @�  B  A�  @@  A�  BH  A�  D0� C?  Dv� Eo  Ap  AP  ?�  @�  B  AP  Bh  Bt  @�  @�  @�  @@  A�  A0  D  A   B�  A�  @@  @@  AP  A�  BX  A�  A�  A0  ?�  @   @�  @@  @�  @   A0  A�  B4  A�  @@  @�  @   @   ?�  B  A�  @@  @   ?�  A�  @�  A�  A�  A@  A`  C�� C̀ C  BL  D@ C�� B�  Ei� L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       123L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       u=�T���Lg?7(|B{|«X9�ѰyA��C=����A�{���@?�E��v^A��B��[Ca���\Z�B� ��&�zаB6��A�Ɏ�B��?�\B>1��ނ�J�x���BVB��¸z�>�` C�4�A��@��;PC�G B o�3���^�F���Bp�B�Z�R��j��O>=�B���B����{t#B;���b��Bۧ�BS5Y�C2�jA�	C��`B���B��K�蠇A�R��g����B�"��4A]���%U��/�fB�IM��S4�U��B#�@��a�u��0KA�qA��:�ƍ�@�RB7|�As����OA���R�4?���rC BA3��aA�qh��x�f[}A$`�B�Aa���?yz����G.@�BB��B���SO2�����1��ծB�
?��Bt�Cd��/�'BxJ�A#,YA��!@� ��*4�$=�L       
categories[$l#L       >                             
                      	                                                      	   
                           	                                           	   
            L       categories_nodes[$l#L                	   
               $   3   6   ;L       categories_segments[$L#L                                                                       &       '       ,       0L       categories_sizes[$L#L                     
                                                                      L       default_left[$U#L       u                                                                                                  L       idiJL       left_children[$l#L       u               	                                    !   #   %����   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K����   M   O   Q����   S   U   W   Y   [   ]   _   a   c   e   g   i   k   m   o   q   s��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       uGҵ�I$V;H$@tH�k
H�>H:�VHE-H��HÈ7H*�uI	�8H+�0HmoH���I� H���G8;EH{�H�d    H	%�G�a^H�� H.�_H�/>H�F�IQ�H�мH���I��G��Fԩ�H?�E,|E9�H�'�H:��HY�lG��q    G�bGC�GC~    H8,H>'=H�_ H̥gGԲ:H���H|]^I/ H�M�H?
~H���H췄H���H�b�H`�2D���F�~                                                                                                                                                                                                                                L       parents[$l#L       u���                                                           	   	   
   
                                                                                                                                   !   !   "   "   #   #   $   $   %   %   &   &   (   (   )   )   *   *   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <L       right_children[$l#L       u               
                                     "   $   &����   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L����   N   P   R����   T   V   X   Z   \   ^   `   b   d   f   h   j   l   n   p   r   t��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       u@      ?;�m   >��?o@�  @�ff>H�9      >��H   ?z�?���>��D��    ?L�D�zа=�
=>�hs=49X@�v�   >P�`?S�F>�I�?|�   D�� BR  D�  D�� B  B8Q�   >�ffB�  ���B��{>D��?ȴ��j=���?�>%=� �@�  B�33?+�   E}  @@     D�@ @@  B�
=>s�F   A�  A�R��g����B�"��4A]���%U��/�fB�IM��S4�U��B#�@��a�u��0KA�qA��:�ƍ�@�RB7|�As����OA���R�4?���rC BA3��aA�qh��x�f[}A$`�B�Aa���?yz����G.@�BB��B���SO2�����1��ծB�
?��Bt�Cd��/�'BxJ�A#,YA��!@� ��*4�$=�L       split_indices[$l#L       u                                                  
         
                                
                            
                          	   	                                      	                                                                                                                                                                                                                                       L       
split_type[$U#L       u                                                                                                         L       sum_hessian[$d#L       uE�8 C0  E׸ B�  B�  E� C�  A�  B�  A�  Bp  E�� D@ C�  B�  A�  @�  A�  B  @   A�  A�  B,  E� B�  C�  C!  B�  C#  BT  A�  @�  A@  @@  @@  @�  A�  A`  A�  ?�  A�  A  A   @@  B   E�  B  Bp  A�  B�  C�� C  A�  A�  B�  Ap  C  A   B4  @   Ap  @@  @   ?�  A0  ?�  @   ?�  @   @@  @   A`  A0  @�  A   A   A0  A�  @@  @�  @�  @   @�  @   B  E�� C�  @   B   @@  Bd  A�  @�  B�  @   B�  CB  B�  B,  AP  @�  A�  A@  B@  A�  @�  A   C  A�  @�  ?�  A  B  ?�  ?�  @@  A@  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       117L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       K=��y��u�A��u���Bl������B�i�dv?��B0��y�BC��B?�z��i�A��@bnV�dE5A���B�m�B殲��J�B�/O��g�?Ц��<�@�G:C�)2@#��B�9DB��=���&B�^���BFt`B��w�iA�rCF��B�I
B���W@�g>�-��A�&����A������w�Cd(��Z?��B1����3A~̮C3#��/��q��.��B�AfU+�fG�A��w@zf¬"���p�ƫA��@?U��B�M�B&�>�o!B2;'����´=���T�L       
categories[$l#L                                                                                L       categories_nodes[$l#L       	         
               #   'L       categories_segments[$L#L       	                                                                L       categories_sizes[$L#L       	                                                               L       default_left[$U#L       K                                                             L       idiKL       left_children[$l#L       K            ����   	               ����                  ����   !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =����   ?   A   C   E   G   I����������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       KG��G��PH4f�G�O    HE�qH�KuH�BPHIQ�H�cuH�N�    H�i�H�b�I�J�H�s*H���G�y    GIXRH*ǆG��HkrH���I',�H�5?J%[H���I8I9�LHʺXF���G�OE~��    HsGt��G��GʝFz�G��                                                                                                                                        L       parents[$l#L       K���                                                     	   	   
   
                                                                                                                             !   !   #   #   $   $   %   %   &   &   '   '   (   (L       right_children[$l#L       K            ����   
               ����                   ����   "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >����   @   B   D   F   H   J����������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       K?� �@��Bt     Bl��   B|  ?p�A   @�   C��   BM�A�  A   =��w@��RB�m�B@�D��    @@  D��    >�b@�  >��   A0  BT  @   D�� @?
=B��w   @�  @@  D�`    B�  @�g>�-��A�&����A������w�Cd(��Z?��B1����3A~̮C3#��/��q��.��B�AfU+�fG�A��w@zf¬"���p�ƫA��@?U��B�M�B&�>�o!B2;'����´=���T�L       split_indices[$l#L       K                                                       
                                   
                                                                                                                                                                                 L       
split_type[$U#L       K                                                                  L       sum_hessian[$d#L       KE�8 E٠ B�  Eِ @   B�  B4  D�� E�� B  B   @   B,  De@ Ch  E�` D:@ B  ?�  @�  A�  A�  AP  D  C�� C[  AP  E�� BL  A�  D4� A  A�  @�  ?�  A�  A   A  A�  @   A0  Cʀ C  B�  C�  B�  B�  A   @�  C�  E�X B(  A  A�  @   C�  C�� ?�  A   A0  A�  @@  @   @�  AP  @@  @�  @   @�  A0  A   ?�  ?�  @   A  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       75L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       W>6T����?0��z-���@@��G�8�_�+4��̬�?��B��@�!|�z<�B| ���wB�a���%?��që�:A�q�C:z����@�t��L2�3BE�BC�\�N����~�A���@��4�);��R^�Ђ�@�i�a �P
B���A?��A�ٵC����A��B1y@[hp��$�B!���v؜��A��h;����͂@9'�f���Vl<�JA����xU?j_A�4�6��ARr�B��9A�-A�Ǵ��A����-�HB9�hC�9B{��J��A(�B<~�AM�K¯?�@�v���?�������j@�L_Cc��]�B�o�m�UB
QhL       
categories[$l#L       $                                      	   
                                         	   
                             L       categories_nodes[$l#L       	                     !   #   &L       categories_segments[$L#L       	                                                  !       "       #L       categories_sizes[$L#L       	                                                               L       default_left[$U#L       W                                                                      L       idiLL       left_children[$l#L       W         ����      	                                    !   #   %   '   )   +   -   /   1����   3   5��������   7����   9   ;   =����   ?   A   C   E   G   I   K   M   O   Q   S   U��������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       WG��GɲG�d�    G�e�H��$H�MTG��H	�xIKI��H���I�GAt�G��[D��Fi� H��(IoBI��ILH��H���I
jI]��G	2v    G�M�G�"*        E���    I>גI9aGT�    H�I<zHL3I�ɋH�+�H���I ��H�͔I��I���I��IHd�                                                                                                                                                        L       parents[$l#L       W���                                                     	   	   
   
                                                                                                               !   !   "   "   #   #   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0L       right_children[$l#L       W         ����      
                                     "   $   &   (   *   ,   .   0   2����   4   6��������   8����   :   <   >����   @   B   D   F   H   J   L   N   P   R   T   V��������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       WA�  =� �>(���z-   @�Q�Ap  =�^5   @�ff>!��=�S�@���D�� D��       Ap  BV  @�A (�>���>A�7@�G�@�     BC�\B�     A���@��4@�  �R^   >�u   �P
>I�^   ?�7Bt  D�  @D�B̊=D�@ A   A�  D�� ?���A��h;����͂@9'�f���Vl<�JA����xU?j_A�4�6��ARr�B��9A�-A�Ǵ��A����-�HB9�hC�9B{��J��A(�B<~�AM�K¯?�@�v���?�������j@�L_Cc��]�B�o�m�UB
QhL       split_indices[$l#L       W      
                                                                                                                                                        
                                                                                                                                                        L       
split_type[$U#L       W                                                                              L       sum_hessian[$d#L       WE�8 C  E�� @   C  EG� Ei� B�  A`  E1� C�  E� D�� A�  B�  @@  A0  E1P @�  C�� A�  C3  E
� D�� CF  Ap  @@  B�  A0  @   ?�  A  @   C�  EP @�  @   B@  C�� A0  A@  B�  B�  C�� D�@ Dm  CC  C   B�  @�  A   B�  AP  @�  @�  A   ?�  C�  B�  E	 C  @   @   Ap  B  C  C  A   @@  A   @   @�  B�  Bp  A@  C�  @�  D>� D�� D@@ C3  C=  @�  B�  B<  Bt  A  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       87L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       i>C�AR"��9j����A�x�9�?i���I�B��C��A���C)����$A���׿$A`������̎�C
M&Br/CC`�����A�̓�RT�C`*����aK��o�B�E�®r��T�,@D��C�/B�L~�&��13�@���Cw�=Bk��B,[��|�@���BćBC'iz�J5�A��iC�\T��f���!� wAE��[�C�G�A��C �]�?����x�C	�鿱��A� ���=�o�B�Z$@dt�n��B�wD���gAɜ8=ögA�rT��g���a½V�A%Tl�!�AY�B�=D�#��B��_��igB-���'��C%��A��@ y���}6@x�B������Bsr|C.�AY����9�B��C'A�:���>B	���{>�K���Q AB�rپ���B{f!L       
categories[$l#L       )                  	                                      
                   
                                        	   
         L       categories_nodes[$l#L             !   "   &   .   1   4L       categories_segments[$L#L                                           	              L       categories_sizes[$L#L                                                        L       default_left[$U#L       i                                                                                                L       idiML       left_children[$l#L       i               	                                    !   #   %��������   '   )   +   -   /   1   3   5   7   9   ;����   =   ?��������   A   C   E   G   I   K   M   O   Q   S��������   U   W   Y   [   ]   _   a   c   e   g����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       iG�8H���G�DH���I���IN'H��yH���H*�cH��,H��I �IX�I7��H�jH���I#F��&G��        H���H�K�H�T�I4�G��0H�3�IN[�I-�PI�AH���Hv�    H{Hw�        G��Fe5�F�P.Gn `IK��IR��G��G)<hHf VH͑�        I�I'�IM�AI<�I���I'ޒI�BILY�IjӬHY^{                                                                                                                                                                                        L       parents[$l#L       i���                                                           	   	   
   
                                                                                                                     !   !   "   "   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   :   :L       right_children[$l#L       i               
                                     "   $   &��������   (   *   ,   .   0   2   4   6   8   :   <����   >   @��������   B   D   F   H   J   L   N   P   R   T��������   V   X   Z   \   ^   `   b   d   f   h����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       i=�hsD� >+B�  D�� D�` >-VBDp�=��?.{>?|�>bND��    >0 �@@  >/�C  >/�Br/CC`��=T��=u<ě�>��B  ?�&�B�  >`A�B�  >1&�B
ffC�/      �13�@���B�     BF  =�\)B�33B�  @   @�  =�
=   ��f���!   B�  B�     >��h=�x�>�x�>#�
@�  A�  A� ���=�o�B�Z$@dt�n��B�wD���gAɜ8=ögA�rT��g���a½V�A%Tl�!�AY�B�=D�#��B��_��igB-���'��C%��A��@ y���}6@x�B������Bsr|C.�AY����9�B��C'A�:���>B	���{>�K���Q AB�rپ���B{f!L       split_indices[$l#L       i                           	         	                                                                                             	                                                                                                                                                                                                                                                   L       
split_type[$U#L       i                                                                                                  L       sum_hessian[$d#L       iE�8 C�  E�x C  C�  DY� E�H C  A�  @�  C�  A�  DR@ D1@ E�  B�  B\  @@  A`  @�  @   AP  C�� A   A�  @�  DQ@ C� Cn  BD  E�� B�  ?�  A@  B,  @   ?�  @�  A  @�  A   CL  B�  @�  @�  A   A  ?�  @@  C�  C�� C�  @�  C
  B�  B   A  A�  E�  A�  Bh  @�  @�  @�  B  @�  ?�  @�  @@  @@  @   @@  @�  C*  B  B`  A0  ?�  @@  @�  @   @�  @�  @�  @@  CC  C�� C�� @�  C߀ A�  @@  @�  C  A  @�  B�  A�  A�  @   @�  @�  AP  E�� @�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       105L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       w>`N�@�v� o���A������?��@�uJ��oA��Cq�P�["<�"(�Bͫ�>�&T��{�B�Vu?oV�³q�D��B �D�5&rD1eTA�(k��k�����Cm����]7A��R���@�n�Bs��C��,A�п�C�����)c�A�y�p��,Bj���i�A��B���C���@��>C#�AS]v ��%���K�!�.�Bn�C���A�ϹA܀�FBB^���%��I�������I�N�\@&8���h@�@�C	��A��P�.2g�Yx��+��fZ�AW��@��2�q�f��A�Ӭ@ ���j��@(C2���0A�3�3�W��$�YH�A�T����B��g�@��CA��AC�����<A'���:@ih�@�� �uU �����`TA����@f���3C��B�]�����B��2��1� 7A�V
������n�@g����O��t�A�}�Y��L       
categories[$l#L       *             
                       	   
                               	   
                                                      
      L       categories_nodes[$l#L                         %   +   ,   3   6   ;L       categories_segments[$L#L                                                                                     !L       categories_sizes[$L#L                                                                                    	L       default_left[$U#L       w                                                                                                      L       idiNL       left_children[$l#L       w               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C����   E   G   I   K   M   O   Q   S   U   W��������   Y   [   ]   _   a����   c   e   g   i   k   m   o   q   s   u��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       wG��H�RPH�"GI *�I�I<ͼH�hvH��Ib��H��,I��I�I3��IW0�H���H�I��$H���I��tII5IIPe8G�L�H�-�I$QFIQӠH���H���I��H�II�HΟ�H�?)H�mI��    H�I�H��IE�sI�?�H���I��H�,�IM��F4�F�B�        IC/gI���H�ӒIX��G/��    H�"�H��H���H"��G��6GV�HI �I.�dIm H��[                                                                                                                                                                                                                                L       parents[$l#L       w���                                                           	   	   
   
                                                                                                                                         !   !   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   /   /   0   0   1   1   2   2   3   3   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <   =   =   >   >L       right_children[$l#L       w               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D����   F   H   J   L   N   P   R   T   V   X��������   Z   \   ^   `   b����   d   f   h   j   l   n   p   r   t   v��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       w>ٙ�@B�\?	x�@�>׍PA@  ?
~�?��   @   >���   AP  D�� =�`B=��D�� @�  >`A�Bb  B7��=��B@�A     >�RA     B  >hs>O�   ?;"�@�  C��,>�D�     =�\)>�t�D�  B.  ?�A�      B���C���=y�#A   ='�?���   �K�!>�ƨ   D�� @@  A`  D�     >-V>	7L>n���I�N�\@&8���h@�@�C	��A��P�.2g�Yx��+��fZ�AW��@��2�q�f��A�Ӭ@ ���j��@(C2���0A�3�3�W��$�YH�A�T����B��g�@��CA��AC�����<A'���:@ih�@�� �uU �����`TA����@f���3C��B�]�����B��2��1� 7A�V
������n�@g����O��t�A�}�Y��L       split_indices[$l#L       w   
      
      
      
                                     	                                                                                                                                                                                                                                                                                                                                                                              L       
split_type[$U#L       w                                                                                                            L       sum_hessian[$d#L       wE�8 E.0 E�  D�� D�� D4@ E_0 D�� C�  D�  A@  D+@ B  A�  E]P D�� B�  C�  C:  C�� D?� A   @�  C�  Cǀ A   A�  A�  A@  DI� E*� B�  D�  B�  ?�  CT  B�  B�  B�  C\  C  C�  C�  @@  @�  @   @   C�� A�  C1  C^  @�  @@  Ap  AP  A   A   @�  @�  C�� D@ C;  E@ B�  A�  Dz� A�  Bl  @�  C  B�  A�  BH  A�  B�  A�  B�  C
  B�  B�  BT  Cw  BD  C�� C  ?�  @   @�  ?�  A�  Cq  @�  A�  A�  C  C  B�  ?�  @�  A  @�  A  @�  @   A   @   @�  @@  @@  @   @�  C(  B�  B�  C� C  B  B@  E@ L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       119L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       q>K�j���rA���z���� ��A��Y�X�?���0�F�zd��*������B��$A3x'��CM�{@P�>���] Ö=	C�E��S�@�����[B���߭�C��B�v�B�p��p��}�����B��hAl.�?�j�B�,�AcR���KC����J��á��A���C�b�L�MÃ �B+FL��`�±��y�F�5��h��C`��B�V�CPQB3��A�TC4]��;��B��K��_AQ���	��ſj�@�j�BK���l�AXd��b���M�@'x$�">gB������<���������%t����eA �>F����PzB;���BZ��A�9�ǆ�'����A-���� @�`M���;���m�¢�B:�BjЗ°6�@Nl�B�������A�����5�Ba�$C�SAݦW����@�n�@q��B�@�L       
categories[$l#L       (                                                                    
                                         	   
               L       categories_nodes[$l#L          	   
                  $   (   *   +   2L       categories_segments[$L#L                                    	       
                                                 'L       categories_sizes[$L#L                                                               	                            L       default_left[$U#L       q                                                                                                    L       idiOL       left_children[$l#L       q               	                                    !   #   %   '   )   +   -   /   1����   3   5   7   9   ;   =   ?��������   A   C   E   G   I   K   M   O   Q����   S   U   W   Y   [   ]   _   a����   c   e   g   i   k   m   o����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       qG�vI�H��IHO �I�H�{(IC��HJ��H �%I ��I=��H�SH�fI���H��H'<�FCa�H�T?I;�H��G� IKnaHˢ`H�vjG��H    H�?�I��H[��HʘH�6SH71�Hi�.        H[C�H��H�\I?6�G�G�kHD �PG1��C�U    H�͚H���Ii�H�YwGX��G�j�G��H���    H�E�H��CH(��H��uI'�H���H��}                                                                                                                                                                                                                L       parents[$l#L       q���                                                           	   	   
   
                                                                                                                                   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <L       right_children[$l#L       q               
                                     "   $   &   (   *   ,   .   0   2����   4   6   8   :   <   >   @��������   B   D   F   H   J   L   N   P   R����   T   V   X   Z   \   ^   `   b����   d   f   h   j   l   n   p����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       q?@  ?;"�@�\)@   ?˅A0  @��RA0  @��      @;dZD�@ >�ff?Qhs      @�(�   D�  =ȴ9BH��B�  @   @�  B��   =�Q�   >�5?B̊=D�� @�  B��hAl.�>�$�   >\(�@�(�@8��   B        C�b@@  ?)��B�  >O�B\)   >�A�C  C`��B�  B(G�>���D�� >�z�>ڟ�?z���_AQ���	��ſj�@�j�BK���l�AXd��b���M�@'x$�">gB������<���������%t����eA �>F����PzB;���BZ��A�9�ǆ�'����A-���� @�`M���;���m�¢�B:�BjЗ°6�@Nl�B�������A�����5�Ba�$C�SAݦW����@�n�@q��B�@�L       split_indices[$l#L       q                                           
                      
                                                                                                                            	      	                                                                                                                                                                                                                L       
split_type[$U#L       q                                                                                                     L       sum_hessian[$d#L       qE�8 E�@ D�� E�� B�  D� C�  B�  E�X B  BT  D  B,  B�  Cπ B�  @   E�� D�@ Ap  A�  @�  BD  C�  A�  ?�  B(  A   B�  Bx  C�� B  B  ?�  ?�  E�P B�  D	� D%  @�  A  @   A�  @@  ?�  B(  @�  C+  C�� A�  @@  A�  A`  @�  @�  A  Bx  B  A�  C�� A�  A   A�  A�  A   EX� D�� B�  B  C{  C�� C�� C�� @@  @@  @�  @�  ?�  ?�  @@  AP  @   ?�  B  A   @�  ?�  C%  @�  A�  C�  @@  A�  ?�  @   @�  A�  AP  ?�  @�  ?�  @�  @�  AP  BD  A�  A   @�  A�  B�  CM  A�  @�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       113L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       u>R|@��j���A��V�w֧�^2?S��@sF�B����ȝB*5����lB]c�Bܦ�>��!xnA��"B�C$��&�<C����$�C(��C��2�ԨLC�dz���wC��i�#o�?�"���%B�0��B2¤r�BO����C�
B��kA�_��DD�}A	G ��"�Bi>CzY�B���B�@�� ��B@�q��DC���¬��¤bC�(�B�m3C���B�z¡澊X�B6ͼð�`��}&�G�B�NA�`�1�_��l�A�J���oA�biB��@����g�;jC���k~g����B�;V@@S�B�qd���@�WSgC����S��Bg0�A���o�ZA��&��6��!@2B���B�J@g��?W|AێA�2�C6	����g!C
G�@+Q�B'��N�B���A�i�� ��B<G�>Hs���R��X@A��A��Z�gbA"I��{L       
categories[$l#L                           
               
                                      	   
                    L       categories_nodes[$l#L       	             +   1   7   8   <   >L       categories_segments[$L#L       	                                                                L       categories_sizes[$L#L       	                                                               L       default_left[$U#L       u                                                                                                        L       idiPL       left_children[$l#L       u               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y����   [��������   ]   _   a����   c   e   g   i   k����   m   o   q   s������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       uG�s�H�a>I#pIH�I˚Iu�`H��H�I�:I�III��Ij�I��EH�VOHB��I�;IK��I�h|I�T�I0%�I���I%�I`��H#AI0�nIg�8I_�H"�H� BH�]�I��IL�Ie�I(�H���I�Hs��I�S:I�9I1�IH��JI I�H�e�H/X(    Iٜ        Hu�I/��I���    H�H:<G�F�� G��S    H�qIs��I-=BH��m                                                                                                                                                                                                                        L       parents[$l#L       u���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   .   .   1   1   2   2   3   3   5   5   6   6   7   7   8   8   9   9   ;   ;   <   <   =   =   >   >L       right_children[$l#L       u               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X   Z����   \��������   ^   `   b����   d   f   h   j   l����   n   p   r   t������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       u>��>bN>�n�>Z�>��P@�  >�t�D�  =�1>��\A�  <�9X@�Q�>�oB�  >�?˅=���>\)?�=q   >�1'@      >oBt  @D�>$�A�  B�Ǯ>�9XA      >#�
@�  >^5?B�  >�dZ>�V?��
>�(�B  @�     ?%�CzY�D�� B�@�� ��   A  D�  ¬��>�1@_�w      @   ¡�B�     =�Q�   �G�B�NA�`�1�_��l�A�J���oA�biB��@����g�;jC���k~g����B�;V@@S�B�qd���@�WSgC����S��Bg0�A���o�ZA��&��6��!@2B���B�J@g��?W|AێA�2�C6	����g!C
G�@+Q�B'��N�B���A�i�� ��B<G�>Hs���R��X@A��A��Z�gbA"I��{L       split_indices[$l#L       u   
      
   
         
         
                  
                            	                  
                
               	             	                                                                                                                                                                                                                                                                                     L       
split_type[$U#L       u                                                                                                            L       sum_hessian[$d#L       uE�8 D�@ E�� DL� D  CZ  E� D@ C=  Cˀ C  C  Bl  A�  E�P C5  C�  B�  B�  CÀ A�  B�  B  @@  C  A�  B(  A   Ap  E�� C  Bh  B�  C�� B�  B�  @@  A�  BL  B�  C�� @   A`  B  Bh  ?�  B  @   ?�  A�  C  Ap  @   B  @�  @�  @�  A@  @@  E� C6  A@  C  B@  A   BD  B�  C  Ci  BL  A`  A`  B�  ?�  @   Ap  A   A�  A�  B�  @@  CK  B�  ?�  ?�  @�  @�  AP  A�  BL  @�  A`  A�  @   A�  B�  A@  A   @�  @   B  @@  ?�  @@  ?�  @�  ?�  @�  @�  E�� B�  B�  B�  @@  A  B�  B$  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       117L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       q>���@0&�����>U�_BZ�����r��ϫ1A��A���C ��ÂEB�>bA&���6�m�[$"�D��@���B�3B�������DC�
�A��������[B��j?��C ���k�������.@���ú3#�B����K
A�SC��b��(]Cerw�XL�B��;B��fæ�lD��B��QBE�M��$����Tt¾\�BѪ�.#�A���B;�C�������W@�����>@���{k:?�5�B_�1�8�<�\�A�zLDBC���v���1��,oA���¬��B�\��#�;�'|��A\AL�B��k��"7A)��BE����F®~�B����\���
�C*�B�� B��S���A�ɝ@e���8�4�	  @r?��A�gK�Ti�B���m�BM7qC?��@�ƞ��*�@��g�l[���1[@� ��?��%��L       
categories[$l#L       &               	                                                                                                
         L       categories_nodes[$l#L       
   	                     #   /   6L       categories_segments[$L#L       
                             
                                          L       categories_sizes[$L#L       
                                                                      L       default_left[$U#L       q                                                                                               L       idiQL       left_children[$l#L       q               	                                    !   #   %   '   )   +   -   /   1   3����   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]������������   _����   a   c   e   g   i   k   m   o����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       qG���I�*H��Hb~�I[�I0� HhJHI�AI��I0hJ��In�Hd�Iz��H�j�HNC�H�h�I1I���I~�9H���I}02I��F�q�Gg�`G�w*    H�8�Iu��H��<H�X�H���I1hG�_�H��bID�H�$�I��I_LH�ɴH��PH�c�H2�IWo�H�(I�pI��D��            Eہ�    I4�tI%��I.��I)|rH���H�dH�mIh�r                                                                                                                                                                                                                L       parents[$l#L       q���                                                           	   	   
   
                                                                                                                                   !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   3   3   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <L       right_children[$l#L       q               
                                     "   $   &   (   *   ,   .   0   2   4����   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^������������   `����   b   d   f   h   j   l   n   p����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       q>�n�>�+>�t�>���B|  ?H1'>��>�E�@�     >aG�   Bb  >�=q>�=qA�  D�� >I�@���?E`B?	�^   ?���   >�/   B��j      >o��@�  ?
��@��@@  >�Q�   A�  ?�T?�9XBx  B�\D�� @��H@   >�\)@�  >�b   ��$����TtB"��BѪ@�z�   >��/Bf  ?�n�D�` >��Bf  @���{k:?�5�B_�1�8�<�\�A�zLDBC���v���1��,oA���¬��B�\��#�;�'|��A\AL�B��k��"7A)��BE����F®~�B����\���
�C*�B�� B��S���A�ɝ@e���8�4�	  @r?��A�gK�Ti�B���m�BM7qC?��@�ƞ��*�@��g�l[���1[@� ��?��%��L       split_indices[$l#L       q                  
   	             	          	                  
                                                	         	   
                                                                     	                                                                                                                                                                                                                   L       
split_type[$U#L       q                                                                                                       L       sum_hessian[$d#L       qE�8 E�  E
0 E� Cc  A�  E� E�� C�� C)  Bh  A`  A   D?� D�� E�p A�  Ck  B`  B|  B�  A�  B  @�  A  @�  @@  D5  B(  C  D�@ E  D�� @�  A   B(  CA  B  A�  B  A�  B�  A�  A   A   A�  A�  @�  ?�  @�  @�  @�  ?�  C;  D@ A�  A`  B�  B  Dq� C�� C� D�� D� A�  @@  @@  @�  @�  B  @�  C,  A�  B  @�  Ap  @   B  ?�  @�  A�  Bp  A�  A   A0  @@  @�  @�  @�  @�  A  A`  A   @@  ?�  ?�  @@  B�  B�  CP  C�� @�  A�  A  @�  Bd  BT  A@  A�  A�  Dj� Cl  B�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       113L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       w>Z�w��@����ТU=BB?�U@�x-� ٢A������C�  B;B+���&��A�X��	�A��@����C���8g�~9�D��¤@PB�Ƿ��H0A�lvCD�g��Y�V=2BE}?�N�A��E�G�U���B�愿�IT�"�A��i�CQ�M����Ì��BY�-�ط�CgR�@Ug�)��A�f��ߛ�B�G�B4�P�/�0}�B���Aߦ�C�l��O��Öd�!.{B���@J��B0�@K]���6A3^��i�P� ��@Z�AA����3@��-�YB$�|�r#�@\����4?�&�I�BX��ň ��3��V4B�[A����g���A���g�w��³������B���&�&]��MG��B"��@��\*�A��)��T@�4��QAQB,<�@}Z0���DB3�$C�A.��?��Ay2���!���)��Rw�Bx����B8�L       
categories[$l#L       (                                  	                        	                                        	   
                        L       categories_nodes[$l#L       	               (   +   .   1   <L       categories_segments[$L#L       	                                    #       $       %       &       'L       categories_sizes[$L#L       	                     	                                          L       default_left[$U#L       w                                                                                                         L       idiRL       left_children[$l#L       w               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y����   [��������   ]����   _   a   c   e   g   i   k   m   o   q   s   u��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       wG��H���H��Hf��HÊ>I4G.H��nHbx�H�f�H��Hr��Iq6�H�ǣIH�7qH��H��pI�I�!HW�(H�G ��HI��H߹4G�z7H�9lH�Z+H��JH�J�H�͙H�I'Ih�H�p�I��H�[<H�3�I`�I/;dIO�GM0�HE�G]X�FQ�E#�F��     G��        FH`�    H<�7H�ARH�XHZ�.H�l�H���H4qmHۥ�H�H]F�b H���HE:                                                                                                                                                                                                                                L       parents[$l#L       w���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   .   .   1   1   3   3   4   4   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <   =   =   >   >L       right_children[$l#L       w               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X   Z����   \��������   ^����   `   b   d   f   h   j   l   n   p   r   t   v��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       w?ļj?��?�n�B>ff   =��w=��-@@     @@  >dZBt  ?	�^=�hs=�{   >���D�� ?St�>���?49X>hr�>bN   B�  >V@�  @@  D�@ B�  Ap  @�  @�  >�Q�??|�=��
?�;BT  @�  >o��   =��wB\)   A�  BY�-   CgR�@Ug   A�f�=�?�-?�+?N�@�\)A�  @�  @@  B4(�   B  =�F@J��B0�@K]���6A3^��i�P� ��@Z�AA����3@��-�YB$�|�r#�@\����4?�&�I�BX��ň ��3��V4B�[A����g���A���g�w��³������B���&�&]��MG��B"��@��\*�A��)��T@�4��QAQB,<�@}Z0���DB3�$C�A.��?��Ay2���!���)��Rw�Bx����B8�L       split_indices[$l#L       w                   	                                   
            	      	          
                                                	                                      
                                                                                                                                                                                                                                                               L       
split_type[$U#L       w                                                                                                              L       sum_hessian[$d#L       wE�8 E�x E� E�� BT  CA  D�� E` E @ A�  A�  @�  C:  C0  D�� Dc� D�� DH  D܀ A@  AP  A@  A�  @�  @@  B�  B�  C  A�  A�  D�  C�� D� C�  Di� D'� C  D�� D%� @�  @�  A  @�  @   A   @   A`  @@  ?�  @   ?�  A   B�  B  B,  B�  B�  A   A@  A�  @�  D�  A�  CR  B�  D@ Bt  C�  B�  C�� C�  B,  D  B@  B�  Cn  DX  C̀ C{  @�  @   @�  @   ?�  A   @   @   ?�  ?�  ?�  A  @�  A  ?�  ?�  @   A   B�  A�  @�  B  A�  A`  B  B  B  BD  @�  @�  A   @�  A@  AP  @   @@  D�� A   @�  A�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       119L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       k>��� ?��,�I��BS[B�3\?�aC@me������
B���@�MC)#�@@�Y�z1CI,��h�A��2Es�Z	���C0d�BC�4�?2�C5���b@C��M@ �|B�Ux�	;_@��B���A�-A D���kA#�C�mH�z¶�A ��0z>�vg�ʈWC��B#"�B�-]����B�}�����@B�$�A`?���nB�>B:; �F̻A,�.JCr�WA�>��[oyB�����^�@�W�hn���Â�����AwƮ@CS9AI�>�7� �"����B�CB	Y����gB!o7@�ʆB�!�A+S-�s�B''�Rg�g�� �T��_�A,ʹ@����Y�?�@���I<���A/��8�A�u�Bެ�B8���[�Adfs@g���}�B8���U�@�j��t|L       
categories[$l#L       $                                    
                                                                	   
             L       categories_nodes[$l#L                
         /   0   1   3   7   :   >L       categories_segments[$L#L                                                                                            #L       categories_sizes[$L#L                                                                                           L       default_left[$U#L       k                                                                                            L       idiSL       left_children[$l#L       k               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =��������   ?   A   C   E   G   I����������������   K   M   O   Q   S   U   W����   Y������������   [   ]   _   a   c   e   g   i��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       kG�1�H�)&H~H���H�#8H;|�Gˁ�H�/^H�d�G�xH:lHC΂H��H}�(H�EgG�4�H���II��H���E��`E��H��>H,�~Hg+�H6&�F��G�АH��I�JH�,HZ�w        H�xI�wMH���I9�H~�I��                G$oPGcF�HS"�HR�F��xG���Fp}    C��l            H��I�HTHa�HE�jH���I	��Hg�#                                                                                                                                                                                L       parents[$l#L       k���                                                           	   	   
   
                                                                                                                           !   !   "   "   #   #   $   $   %   %   &   &   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   3   3   7   7   8   8   9   9   :   :   ;   ;   <   <   =   =   >   >L       right_children[$l#L       k               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >��������   @   B   D   F   H   J����������������   L   N   P   R   T   V   X����   Z������������   \   ^   `   b   d   f   h   j��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       k>$�D�� >1'   >�   ?ǍP<D��=ȴ9A�     @�  ?�z�?�z�>�@E�>%=\Bb  B@  @@     >��>��HB|  @@  ?BJ   @�  >ix�?r�B���A�-@�  B�  >]/BH��=�%=m�hA ��0z>�vg�ʈWA   @�  >)��A�           B�$�   ��nB�>B:;    >��D�     =�S�>>v�?�   @�W�hn���Â�����AwƮ@CS9AI�>�7� �"����B�CB	Y����gB!o7@�ʆB�!�A+S-�s�B''�Rg�g�� �T��_�A,ʹ@����Y�?�@���I<���A/��8�A�u�Bެ�B8���[�Adfs@g���}�B8���U�@�j��t|L       split_indices[$l#L       k   	      	            
                     
   	      	                                        	   	                       	   	                                                                                                                                                                                                                                                                   L       
split_type[$U#L       k                                                                                               L       sum_hessian[$d#L       kE�8 D�@ E�� D{� B�  A�  E�� C�� C�  A  Bh  A�  A0  E�P DS@ @�  C�  B�  Cƀ @�  @�  A�  B(  Ap  @�  @�  @�  E�� A�  C�� D
  @�  @   C� B  B�  @�  C�  B�  @@  ?�  ?�  @�  @�  A  A�  A�  @�  A   @   @   @   @   @   @�  Edp D�` A0  AP  B�  C\  B(  C�  C�� B�  B  ?�  A�  B�  @   @   B@  Cf  A�  B�  @�  @   @�  @@  A`  A  Ap  @�  @�  ?�  @�  @@  ?�  ?�  ?�  ?�  E0  DQ� D\  D� A   @@  @�  A   A  B�  Bx  C  A�  A`  C�� CE  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       107L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       U>m��t�BZV>�����i_�Ҧ�B�@R�I�?�J��v7��B�I:ª��A8CbR}�@0C�?�A��A>Us£I$��4C��>�B���@�#��ac�^~B.W���=�C����7A�Z��)sA��B�d�����B�������?�C�B����[��A8(��B��{®�HAg�����2p�����m�@���C���A����ÓCA��(@����~��-�7?�<B��@'y��F��@���A�Ʊ>n�"�U�A�(����G�(c�Aޫ�?��@-���3 Aa������-A���2����@��A��d����C	:�B�MAv'��KZL       
categories[$l#L       .                                       	   
                                                                                	   
                      L       categories_nodes[$l#L                	                  #   $   ,   2   4L       categories_segments[$L#L                                                                                     *       ,       -L       categories_sizes[$L#L                                                                                                  L       default_left[$U#L       U                                                                       L       idiTL       left_children[$l#L       U               	                                    !   #   %��������   '   )����   +   -   /����   1   3����   5   7��������   9   ;   =   ?��������   A   C   E   G   I   K   M��������   O   Q   S��������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       UG�"G��H6:�Gy�Hu
�H%�_H�l;H�H��EM��H�IYHיG�Y G�rHQ��H���G8I�IF,H/{        HN1�Hc�    GX�F���G"}L    F��Hsu    H���H�K        H��LI��&H֘�H�v        G��xH�F�<Fe�Ek:B�J E���        F߂�G���E�y                                                                                                                                L       parents[$l#L       U���                                                           	   	   
   
                                                                                                           #   #   $   $   %   %   &   &   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   2   2   3   3   4   4L       right_children[$l#L       U               
                                     "   $   &��������   (   *����   ,   .   0����   2   4����   6   8��������   :   <   >   @��������   B   D   F   H   J   L   N��������   P   R   T��������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       U?��m?��   >o��=�-B2  B<=q   >�(�   >.{   @S33   D��    B2  D�� ?}p�£I$��4>�   B���   @�  @�  B.W�@   @n{�7B2  B,  A��B�d�      D�� ?���B����[��@�  BR  B�\   @�  B@�A"�\�����m�   B|     �ÓCA��(@����~��-�7?�<B��@'y��F��@���A�Ʊ>n�"�U�A�(����G�(c�Aޫ�?��@-���3 Aa������-A���2����@��A��d����C	:�B�MAv'��KZL       split_indices[$l#L       U   	                                     
                                                         
                                                                                                                                                                                                               L       
split_type[$U#L       U                                                                        L       sum_hessian[$d#L       UE�8 E�p Bd  E�  B�  A�  A�  D� Eň @�  B�  A   A�  A�  A   D  @@  C�  E� @@  ?�  A   B�  @   A   A   @�  @@  A�  A  ?�  C-  Cπ ?�  @   C  B�  D@ E�@ @�  @@  B4  BT  @�  @@  @�  @�  @@  @�  @�  AP  @�  @@  B�  B�  C  C�� A�  C  B(  B�  C�� C`  B�  E�� A�  A�  B  A�  @@  @   ?�  @   @�  @   @   @   @   ?�  @�  A  @�  @   @   ?�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       85L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       o>�QAXT)�;�A���%���\��^��A��3B�YL�]�BX����P����B��w����B��4��-C]��9��(����i B���Z��C!'�ý�����̰�C�"�A�I���I�Baޏ�l��_LÖ��C�o�혅C��A�(��o��tz'�֏���W���ށA!T@leUBG����Al��C�B<A��pA�.��uB%�[�#s��#�B{ϠB��C�,Cw�A���£8�����A�_!���� �B �s��SA{���噴�Ǚ6A6��B���Ѷ$�W�7Bx>UCC��B-���;�<�����BeV��&~vA~g���g�jUx?������A��_A��gB���-�aB
���1*B�!��ݏ�B#@��B�#M?Μ�A�T>��C��A��A{��P;��|0�� ߴ���=M^L       
categories[$l#L                   	                                  L       categories_nodes[$l#L                         -   1   9L       categories_segments[$L#L                                           
                     L       categories_sizes[$L#L                                                               L       default_left[$U#L       o                                                                                                       L       idiUL       left_children[$l#L       o               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M��������   O   Q��������   S����   U   W   Y   [��������   ]   _   a   c   e   g����   i   k   m������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       oG�H�H��H�6H�O�G�H�̃H;o�IvIH�HNG�D�G!�II_�Hߍ5I��H&�H�#H� �H��xH���E?@G��F�<�F�LH���H�EH�16H��H|z~G�(H��I�I'��IRVG��$G3V GO�\GW�`H�L�G���        G��H\�        E��    H���H��-H��6HJk        G��G��H��oH�XE��fG�V�    H�VI���H��&                                                                                                                                                                                                L       parents[$l#L       o���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   $   $   %   %   &   &   )   )   *   *   -   -   /   /   0   0   1   1   2   2   5   5   6   6   7   7   8   8   9   9   :   :   <   <   =   =   >   >L       right_children[$l#L       o               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N��������   P   R��������   T����   V   X   Z   \��������   ^   `   b   d   f   h����   j   l   n������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       oD�`    D�� ?L�DB�  >�D�@ >["�>M��=��P=���>k�   >�$�?�>ix�BM�@  >��@�  >�u   >���>/�>�   >���?���   D�` ?#�
?C�
>�uD�` =�?aG�=���B�  Bd  �o��tz'B8  > Ĝ��ށA!T   BG�@�  A�     =8Q�A�.��u>��B\)>ٙ�=���   @   Cw�?Z^5@�  D� A�_!���� �B �s��SA{���噴�Ǚ6A6��B���Ѷ$�W�7Bx>UCC��B-���;�<�����BeV��&~vA~g���g�jUx?������A��_A��gB���-�aB
���1*B�!��ݏ�B#@��B�#M?Μ�A�T>��C��A��A{��P;��|0�� ߴ���=M^L       split_indices[$l#L       o             
      	                  	                     	      	      	                                     
                          	                                                	                                                                                                                                                                                                                   L       
split_type[$U#L       o                                                                                                       L       sum_hessian[$d#L       oE�8 Cր E�� C�� B�  C   E�� C�  B  B�  A0  B�  A�  B  E�� C�� A�  A�  A�  @�  B�  @�  @�  B�  A�  @�  A�  A�  @�  Cy  E�� CQ  B�  A@  A0  @�  A  A`  @�  @�  ?�  Ap  Bh  @   @   @   @�  B  B  A0  A0  ?�  @�  A@  AP  A   A�  @   @�  ?�  Cx  B�  E�X C'  B(  BH  A�  A   @�  @   A  @�  @@  @�  @�  A@  @   @@  @�  A  @�  @   B`  ?�  ?�  A�  AP  A�  A�  @�  @�  @�  @�  @�  @�  @�  A   @   @�  @@  A�  ?�  ?�  @�  ?�  Cr  @�  B�  @�  A�  E�p L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       111L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       S=�n�B�s>�d��5h�A^��A��X����LSg@nr��7�KB��BL�"�D*���>�����4��AVz����@�KnB�bvCu�G�@�R�Wé�����0�_��BF�P����B��D�0M@A.�M�H�
C B�_`Cl�'��=�j�Ak8�A<C��(�WU�5¸�
A��"C�z�v4@����2AL9�By$@_?4�����Y �ܱ�@ڠMA��'B/��Cw!����B�e�º��@�uBy����tBbaB��.U»��@����u������f�A����A��A7GB�dA����
 �=˾AZ�
���qA���L       
categories[$l#L                                                L       categories_nodes[$l#L       	      
            !   )   ,   .L       categories_segments[$L#L       	                                           	       
              L       categories_sizes[$L#L       	                                                               L       default_left[$U#L       S                                                                         L       idiVL       left_children[$l#L       S               	         ����                  ��������         !����   #   %   '   )����   +   -   /   1   3��������   5   7   9   ;   =   ?   A   C   E����   G   I   K   M   O   Q����������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       SG���H}�G��(G7lG���H���H���DM�     G�T�H0"II��I
�[Hu�TH��        G8	^G1X�GPN�    I4hH�GH>txH�x    H+�7H�rG��D�3�E��6        D��D���Io�I�DH5L�H��HT:H>�gEMG�    HO�G��I�cHl�*H��H'�                                                                                                                                        L       parents[$l#L       S���                                                     	   	   
   
                                                                                                   !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   +   +   ,   ,   -   -   .   .   /   /   0   0L       right_children[$l#L       S               
         ����                  ��������          "����   $   &   (   *����   ,   .   0   2   4��������   6   8   :   <   >   @   B   D   F����   H   J   L   N   P   R����������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       S<���>0 �=���?49X>n�B  =���   @nr�@@     ?St�@�=��
=�^5���4��D��    >�=qB�bv?'+?�  =�O�B4(����0?���D�  >��`      A.�M�H�
   B33@@  A�  @�  D�� D�  @      �5B�     ?�bN   >�+B�  AL9�By$@_?4�����Y �ܱ�@ڠMA��'B/��Cw!����B�e�º��@�uBy����tBbaB��.U»��@����u������f�A����A��A7GB�dA����
 �=˾AZ�
���qA���L       split_indices[$l#L       S            	                                	                            
                                                                                                                                                                                                                                L       
split_type[$U#L       S                                                                          L       sum_hessian[$d#L       SE�8 A�  E�H A  A�  C<  E�h A   ?�  AP  A   C  BX  B`  EԨ ?�  @�  A   @�  @�  @   BT  B�  BD  @�  @   BX  BX  E�� @@  @�  ?�  @�  @@  @@  B  A�  A   B�  B,  @�  @   @@  B  A�  A�  A�  E�P E	P @   ?�  ?�  @�  ?�  @   ?�  @   A�  A   Ap  @�  @�  @   @�  B�  @�  B  @@  @@  ?�  ?�  B  @�  @�  A0  A�  @�  A`  A�  E�8 CC  E� B0  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       83L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       m=���?�G��?���;A���R�pB�3?%l��N�C/[�A*��C.����HB�mw�O��@��Br��¡CT� � C�d'�b��A��Cd%�AD��A������yBF��P�*�i�C6�����B�b�?�߁C[f�y,�C��KB���¦��C
�B�F$���^@W�UB���.WBB���@������4AT7gB����1�q��{B: �¨�BTL�C+���&C}�tA�6 ��E���+�¤UAm�sBl�q���z@�g�9AB��:��M��5�B�H-A�ûC�/��GF��+�A�z�@6 4�Ě�gB&dA?"MA�X����	�An��¨�GB���|��@w�A&�By_7��}w¬�gBW�IgQ@��
�	�l@���AВ�@J��B����n����>B��I@�E����3A��L       
categories[$l#L       (                                       
               	                                              	   
                       L       categories_nodes[$l#L       
                     '   (   *   8L       categories_segments[$L#L       
                                                         %       &       'L       categories_sizes[$L#L       
                                                                      L       default_left[$U#L       m                                                                                                 L       idiWL       left_children[$l#L       m               	                                    !   #   %   '   )   +   -   /   1   3   5����   7   9   ;   =   ?   A   C   E   G   I   K   M   O����   Q   S   U   W   Y����������������   [����   ]   _   a   c   e   g   i   k������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       mG�_�H�BH�7�H/?�I ˳H�a�HS+�H��IM3�H��NI,ڋG��hH���G�Z�H�H�H��2H=II;$I��{Gs��H��8H�I�=G��E�u=H9ýH�t0    G�gH�u3H0=�H���I;mxH�)}H	7mI���HQO�I[�I��CE�TEzؠ    FC�@H�F�G�kI5T�IN��                G��A    I��Hq��G`_E��DG�(0G��G�PGUh�                                                                                                                                                                                                L       parents[$l#L       m���                                                           	   	   
   
                                                                                                                                   !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   *   *   +   +   ,   ,   -   -   .   .   3   3   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <L       right_children[$l#L       m               
                                     "   $   &   (   *   ,   .   0   2   4   6����   8   :   <   >   @   B   D   F   H   J   L   N   P����   R   T   V   X   Z����������������   \����   ^   `   b   d   f   h   j   l������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       m@�  B�  >���B�  D�    @�  =A�  >�C�D�    >dZD�` >Xb@�  =�         >���B�  D��    D�� >޸R>ՁBF�@@  @�  =�/B�  >��>n�>��A�A  @Q�>t�      C
�   >?|�@   =uD�� B���@������4AT7g>�-�1�q>�C�?X>���   D�  @_\)?&$�>�+��E���+�¤UAm�sBl�q���z@�g�9AB��:��M��5�B�H-A�ûC�/��GF��+�A�z�@6 4�Ě�gB&dA?"MA�X����	�An��¨�GB���|��@w�A&�By_7��}w¬�gBW�IgQ@��
�	�l@���AВ�@J��B����n����>B��I@�E����3A��L       split_indices[$l#L       m                        	                           	                              	                            	                              	                            	                            	                                                                                                                                                                                                L       
split_type[$U#L       m                                                                                                   L       sum_hessian[$d#L       mE�8 E�P C  E�` C�  B�  BX  Eɨ C7  A�  C�  A  B�  A�  A�  D?� E�� B�  B�  @�  AP  A0  C  @�  @�  A�  B�  ?�  A�  A�  Ap  D8@ A�  B  E�� B  A�  A�  B�  @@  @�  @�  A   @�  @�  B�  C1  @�  ?�  @   @   A�  @�  Bh  A@  A�  @�  @�  A  A   @�  D)� Bh  A�  A@  A�  A�  E` EL� A�  A@  A�  ?�  A�  @@  B�  A�  @   ?�  @   @   @�  @@  ?�  @�  ?�  @�  @�  B�  A�  C  A�  @@  B   A�  A  @@  @�  AP  @@  @   @@  @�  @�  @@  A   @   @   @@  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       109L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       m=���AQ�S�87H@���B�K�B�P��M�B*9�����C��?-�!�%�B�\��-L:�L��A��B�\?��±@�CsQCUX��C�m��B����eB��uB����*�_K�>��	�ol�C2�Cm�TA���(�Bqي��fB;E�B��~BJ�HB�	W��?C��BQ-���k����|�E5�B<n+�7`C?/C&a�Èu	�G�A�c�����%�A
P����@�D@P/B���=KgB��vB/���,��ھ��n�B\׷@c���w9���`B~'��LWB&�?[�g@�s�BPL¿{���LBr���>�G4�;�@�:��?4��0gA�bt� 	�A�^�B��B"�Z�?���-\�B�$��8N�����º��d��A)# @���B��4B`$��1^��K�?`03�iC�@��KL       
categories[$l#L                                                                      L       categories_nodes[$l#L                      (   ,   -   0L       categories_segments[$L#L                                                                L       categories_sizes[$L#L                                                               L       default_left[$U#L       m                                                                                                   L       idiXL       left_children[$l#L       m               	                                    !   #   %   '����   )   +   -����   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I����   K   M   O����   Q   S   U����   W   Y   [   ]   _   a   c   e   g   i   k��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       mG�TJH+�G��H�pIE]�H���G�6H���H���I(��H�w2H!�kH�c�H��G�I�H��H��H���H y�    H���H��G�Ʈ    G���H���H�cnH���H��>H��HE�I�NI+�^H`HZ~^H���I'b�G·
    F��#GJ��HtT    G�6�Gc�GM�V    F8Hp�H#�tG$��H��|GV�HK�Hq:�H�??H@-�H�:W                                                                                                                                                                                                        L       parents[$l#L       m���                                                           	   	   
   
                                                                                                                             !   !   "   "   #   #   $   $   %   %   &   &   (   (   )   )   *   *   ,   ,   -   -   .   .   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   :   :L       right_children[$l#L       m               
                                     "   $   &   (����   *   ,   .����   0   2   4   6   8   :   <   >   @   B   D   F   H   J����   L   N   P����   R   T   V����   X   Z   \   ^   `   b   d   f   h   j   l��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       m=�C�=�%=�v�>8Q�D�` B  =��D�� @�  ?^��>w��?�?}=��m@�  >��>)��D�  >���B  >8Q�CUX�>1&�>}�   B��   >�
=BH        A�  =�"�@�  @�  ?U?}D�` ?`BBt  >1'B��~   >$�D�  C��      @�  �E5�   @@  @�  =���B�  B\)@�  ?l�D�  @@  >�M����@�D@P/B���=KgB��vB/���,��ھ��n�B\׷@c���w9���`B~'��LWB&�?[�g@�s�BPL¿{���LBr���>�G4�;�@�:��?4��0gA�bt� 	�A�^�B��B"�Z�?���-\�B�$��8N�����º��d��A)# @���B��4B`$��1^��K�?`03�iC�@��KL       split_indices[$l#L       m                              
      
         
                      	                                               
      	                                                                                                                                                                                                                                                                        L       
split_type[$U#L       m                                                                                                     L       sum_hessian[$d#L       mE�8 C΀ E�P C�  Bd  B�  E�� C  CL  A@  B4  B   B8  BL  E�H B�  B  C  B`  A   @   A�  Ap  A�  @�  @�  B   A�  A�  C�� E�` B�  A�  Ap  A�  B�  B|  B,  AP  @@  @�  A   A�  @   AP  AP  Ap  @�  @   A�  A�  Ap  A0  A   A�  C  C�  E�� D�  B   BX  A@  A   @�  A   @�  Ap  Bd  A�  A�  B8  B   A0  A   @�  @   @�  @�  @@  @�  Ap  @@  A   @@  A   A0  @�  ?�  ?�  @�  A  @�  A�  @@  A@  @�  @�  @   @�  @�  A@  C  @�  A  C�� D�� E%� D  Dp@ L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       109L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       S>#
�A��+��)BR���|µӸ��;xA���CbaA�3�� ϒAx]f�N�6=;N�80s�1O�B�YA{� C�L��?r>B,A��U�]CL B��E�~������e�B�����TcB��CL�BŒ�j�5BtCH�B�2�Bw�m ��_=���\BN�@P?4An��CH�A������J�]@��4�/�KA��UBo:�A��.�k�oA�l�B�57�s�BO��/��$BT��e�B�G?�fB*O�@�G�9��A!8���B����O�iB�j�0� A���BN<tA0�zA�V7�� >�6����A# ��HX����AT6GL       
categories[$l#L                                                   
                                        	   
         L       categories_nodes[$l#L                   $   &   ,L       categories_segments[$L#L                                                  L       categories_sizes[$L#L                                                 L       default_left[$U#L       S                                                                         L       idiYL       left_children[$l#L       S               	                           ����         !   #����   %   '   )   +   -   /����   1   3   5����   7   9   ;��������   =   ?   A   C   E��������   G   I   K������������   M   O����   Q������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       SG|o]H;�*HX��H5^�H�jH�~G��Hk��H�@�H��H,N�G�YeG���G���    HSF�H*6�G�H(�    H��H,��F�5GCRGr�Gi�    G��ZG�5G�9�    G`��H�F��        F.��H�hG�-jHY�pH��2        FY�E��EF�            G�)�HM6Z    F��t                                                                                                                        L       parents[$l#L       S���                                                           	   	   
   
                                                                                                                 !   !   $   $   %   %   &   &   '   '   (   (   +   +   ,   ,   -   -   1   1   2   2   4   4L       right_children[$l#L       S               
                           ����          "   $����   &   (   *   ,   .   0����   2   4   6����   8   :   <��������   >   @   B   D   F��������   H   J   L������������   N   P����   R������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       S=T��>8Q�=]/>p��A�     A�  @�     >KƨB�=qD�� A�  A�  �80s>0 �D�` ?��D�  �?r>B�  BnffA   =�j   B�  ��e?��>��Bt  B��B,  =<j@@  BtCH�   >bN   Bb  @�  BN�@P?4B�33   B
ff����J�]@��4>Ǯ@�  Bo:�A�  �k�oA�l�B�57�s�BO��/��$BT��e�B�G?�fB*O�@�G�9��A!8���B����O�iB�j�0� A���BN<tA0�zA�V7�� >�6����A# ��HX����AT6GL       split_indices[$l#L       S                                                                                                                                                                     	                                                                                                                                  L       
split_type[$U#L       S                                                                             L       sum_hessian[$d#L       SE�8 CY  E�p B�  C   A�  Eՠ B�  A`  Bl  B�  A`  A@  EՐ @   B@  A�  A   @�  @@  B`  B�  @�  A   @�  A  @@  E� A�  B<  ?�  A   A�  @�  @@  @@  @@  BD  @�  B(  A�  @@  ?�  @�  @@  @   @�  @�  @   E�h CU  @@  AP  B  A  A  ?�  A@  @�  ?�  @�  @   ?�  Ap  B  @�  @@  B$  ?�  A�  @�  @�  ?�  @   ?�  ?�  ?�  E�� D�� C'  B8  @   A0  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       83L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       e> ���]��@0:���d��p�B���?Z7��[�R��B,`��v�(¸4BϽ\��8?�>By��2�A���À��B�[a�l�M���B7oA`����{Bn�C��^»��"dBed��3'CX��+¨o�@c=z���g®�_A��SCb���C��C�V�H��A�~By��Âώ�M'B��CsW�A���Cҵ��3N ��C ����C�
�Aް��,��?����sB�W��.��A�3q� ��A�%����A���A��Q����A�h�B����y,#������'<BƄ�?:�n�
��#�A�\�B
��O��A k`��>�)BrB��(Af�{��A���C PDB ���&��A�"z��$M����Bh4C2����|�A�}��겷�~V*A���=���L       
categories[$l#L       +            	                                    	   
                        	                
                            
                 L       categories_nodes[$l#L          	                     )   +   ,   2   3L       categories_segments[$L#L                                                                              (       )       *L       categories_sizes[$L#L                                                                      
                     L       default_left[$U#L       e                                                                                          L       idiZL       left_children[$l#L       e               	                                    !����   #   %   '   )   +   -����   /   1����   3   5   7   9   ;   =   ?��������   A   C   E   G   I   K   M   O����   Q   S   U   W   Y   [����   ]   _   a   c��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       eG�0vH�%LH���H��Hö%I&��HpK�H�	bHu�I�KHk��IP�tI(4SG�.6HV��H�w�H�?�    F.b Ix0H�N�Hl��H��Hڞ�    I �<IQj�    E�N8H���Ha �H���H$e�H��dH���        H��I;��H��LINY�H��]H޷ H�Z�H�~    G�ƧH:�|H��zH�N�G��A�*     H]�IMH��>HX�                                                                                                                                                                                L       parents[$l#L       e���                                                           	   	   
   
                                                                                                                       !   !   "   "   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   .   .   /   /   0   0   1   1   2   2   3   3   5   5   6   6   7   7   8   8L       right_children[$l#L       e               
                                     "����   $   &   (   *   ,   .����   0   2����   4   6   8   :   <   >   @��������   B   D   F   H   J   L   N   P����   R   T   V   X   Z   \����   ^   `   b   d��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       e>z�H<�>�%?^��=0 �=�->8Q�=�F@@     @;dZ>׍PB�  <�/=o   >� �A���B"��>�r�?��   A�  D� ��{      »��   >��=49X   ?�=q@Q�D�  ���g®�_@33>,1A�  =+   >���      �M'B@�?$�/>�=qA         ����Bp  ?�wA   =H�9�sB�W��.��A�3q� ��A�%����A���A��Q����A�h�B����y,#������'<BƄ�?:�n�
��#�A�\�B
��O��A k`��>�)BrB��(Af�{��A���C PDB ���&��A�"z��$M����Bh4C2����|�A�}��겷�~V*A���=���L       split_indices[$l#L       e   	      	   
                                        
                                                                         	                               
                                                                                                                                                                                                            L       
split_type[$U#L       e                                                                                         L       sum_hessian[$d#L       eE�8 E8� E�� Co  E)� B�  Ez� Cg  A   CC  E� A�  B�  A  Ez  A�  CI  ?�  @�  B�  B�  E� B�  A�  @�  B�  A�  @   @�  C#  Eo� A�  A0  B�  B�  @   @�  B|  B  B�  A�  DϠ D?� B�  @�  ?�  A�  A@  B�  A@  @�  @   @�  @�  C  B�  EhP @�  AP  A   @@  B�  A@  B,  B@  B$  A�  A�  Ap  A   B�  A   A  DX� DF� D!  B�  Bt  A�  ?�  @@  @�  A   A   @�  A�  B<  A   @�  @   @�  ?�  ?�  @@  ?�  B<  B�  B�  A0  B  Ee� L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       101L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       q=��+@� ��W�Aj�_�'.��/�,��A��7��݁A,���� �A~��¦-�@ex��?��AsA1C�lÒ{��L��BPX����B��p�*��Bd��}�C�ǳ�ݸ�U�@�5�B�V���TA;�!BǛ5���C� ���z��n����>±4C �A��Ac��«f��ʋ�CG��A�{��v<@��C
�����Z¤PC��A���>�C!�CC��D�Q@�`���X�CCuA濤����A��K@�Y�����As��C��	LBdCA��=���B��:B��)@��@.�[B�����iA���ۉBZ �A�e��ʶB��S��B����
U¢����	@��� ��A��B���Adj��������mw�B���	%e@�m'B�#��^�A��?ψ�A�4��'`z�d��A�#�>��*�ſ�����VAd�ML       
categories[$l#L       H         
                	   
                     	                               	   
                                        	   
                                  	   
                                     	   
                   L       categories_nodes[$l#L                         "   '   ,   -   0   4L       categories_segments[$L#L                                                         ,       8       E       F       GL       categories_sizes[$L#L                                                                                    L       default_left[$U#L       q                                                                                               L       idi[L       left_children[$l#L       q               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E��������   G����   I   K   M   O   Q   S   U   W   Y   [������������   ]   _   a   c   e   g   i����   k   m   o��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       qG�4�H���H`�AI$SH�%�H��2HY�}I�`H�a�H�1 I�vH�3RI���Hh�vH�zH�'IIsQFƯ H?�H���H�XYI(@�I��H�+�D�n Ha;�IE6�H��Hd�H�D�HH=(I��IC��H�/�I/Ō        Ho��    I�=H�w�HW�I�QHR��I5�MI?�H�I@H_H(�            Eu�I%�RH��H�^H/��H�x\H���    H|K�H�v/H��                                                                                                                                                                                                        L       parents[$l#L       q���                                                           	   	   
   
                                                                                                                                         !   !   "   "   %   %   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   4   4   5   5   6   6   7   7   8   8   9   9   :   :   <   <   =   =   >   >L       right_children[$l#L       q               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F��������   H����   J   L   N   P   R   T   V   X   Z   \������������   ^   `   b   d   f   h   j����   l   n   p��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       q>�O�?]/>�>�ZA�        ?Y�D�� D�� D�  ?�@@  A���@@  >���@@     @�  >�bN>E��D�  @   ?��h      D�� D�@ Bճ3>��PA0  >�S�@�  @_\)   ��z��n�A   ±4   >�%?1&�@o�PB!        ?d�/?��   ���Z¤PC��   =�BK��>�z�@�1B�  >�ƨCCuD�` ?�P>�Z@�Y�����As��C��	LBdCA��=���B��:B��)@��@.�[B�����iA���ۉBZ �A�e��ʶB��S��B����
U¢����	@��� ��A��B���Adj��������mw�B���	%e@�m'B�#��^�A��?ψ�A�4��'`z�d��A�#�>��*�ſ�����VAd�ML       split_indices[$l#L       q                                      	                         
                                                                         
                                               
                                                                                                                                                                                                                              L       
split_type[$U#L       q                                                                                                      L       sum_hessian[$d#L       qE�8 E  E�� D�� Dh� CH  E�x D�� B$  C� C� B�  B�  EQ� D�  D�@ B  A  B   C�� C8  BX  Cˀ B�  @�  @�  B�  C  EI� B�  D�� D�@ B@  A�  A�  @   @�  A�  @   A�  C�  B�  B�  A�  A�  B�  C�� B�  A�  ?�  @�  @�  @   B�  A  @�  B�  E>� C.  ?�  B�  D�� B�  D�  B�  B,  @�  @�  A  A  A   A�  @   A   AP  Cj  A�  Bx  BX  Bx  @�  A0  A�  Ap  A   BH  B   A   C�� B�  @   A@  A   ?�  ?�  A�  Bt  @�  @@  @�  @   B�  A   E8� B�  B  C  B   B�  D  C�  A   B�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       113L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       s>(�����p?$m�A�MG�c��weAy�g���sB&]A�	a��1?.����m@�HB`��BC<��`B�;���QBbBk���� @������(@ ��,�A�����$��A$��B����)�?��gA����6�(��u�C]�7B'j�B�
��lIB�@�C%�=A�l�°�Xä	�B=���*�a�K,�A�h�?�/�B:N�B�T�����Ê9���M¯17Bt����)�C4�����B��Tzf����LmB���A�#��.�xB��Ah���P>THB -�S B]I�A,��B
j��Y���4ئ@��M���_��Z?f�{� �{����g�B��T�?(N�#�B�@��2����B�������A
�\@����(o������@�A�WZ�S @��~A��AD���.���/AX�HB�5 �,����"Af,��
gA�mL       
categories[$l#L       d                                
                                                     	   
                                              	   
                                 	   
                                  	   
                                     
                                        	   
                    L       categories_nodes[$l#L                                     $   %   '   4   9   :L       categories_segments[$L#L                                                         "       /       1       <       F       S       a       b       cL       categories_sizes[$L#L                                                                             
                                   L       default_left[$U#L       s                                                                                            L       idi\L       left_children[$l#L       s               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =��������   ?����   A   C   E   G   I����   K   M   O   Q����   S   U   W   Y   [   ]   _   a   c   e����   g   i   k   m   o   q����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       sGv#H��G�3H`
H�"�H�>HrWG��LH��
G��:H���GɁYH���Hh`H�KD��`F��H��G�eHc|VG��EH��Hu�HU�nH`�>H`�HmFG�=�GƃNH��GG]�|        FG�    H��>H5/xDf0�G�HF�b�    E��@GA�-HI��G���    G: 1ISM�I � H�gH��I	��H�ۢHg�H@G(w    G�f�G���G�+uH���G� �Fx�(                                                                                                                                                                                                                L       parents[$l#L       s���                                                           	   	   
   
                                                                                                                           !   !   #   #   $   $   %   %   &   &   '   '   )   )   *   *   +   +   ,   ,   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   9   9   :   :   ;   ;   <   <   =   =   >   >L       right_children[$l#L       s               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >��������   @����   B   D   F   H   J����   L   N   P   R����   T   V   X   Z   \   ^   `   b   d   f����   h   j   l   n   p   r����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       s@      ?;�mD�  >+?)��@�  =���>�7L>Z�?!��A  D�� =�O�      >�bD��    >,1      >n��B�  ?d�/      @@     B�\@D�?��gA���@�
=��u�>7K�      ?�"�   �Bj��=o?�bN@�33B=��@[oBnffB��{?Y�#>Q�D�@    @�p�Bj��D�� ¯17      ?���B�
=D�@ @��\zf����LmB���A�#��.�xB��Ah���P>THB -�S B]I�A,��B
j��Y���4ئ@��M���_��Z?f�{� �{����g�B��T�?(N�#�B�@��2����B�������A
�\@����(o������@�A�WZ�S @��~A��AD���.���/AX�HB�5 �,����"Af,��
gA�mL       split_indices[$l#L       s                        	                                      	                                                        	           
                                                                                                                                                                                                                                                                                            L       
split_type[$U#L       s                                                                                                    L       sum_hessian[$d#L       sE�8 C0  E׸ B�  B�  E�0 C�� AP  B�  A�  Bd  E�� C	  C�� B�  @@  A   B8  A�  A   A�  B  A�  D�  E�h B�  A�  @�  C�  A�  B  ?�  @   @�  @�  A0  B  @�  A�  @�  @@  @�  A�  A�  A   @�  A`  D�  C'  E�� B�  A�  B�  A�  @�  @�  @@  B�  C+  A   A�  A�  @�  @�  @   @   A  A�  A�  @@  ?�  A`  A0  @   @�  @�  ?�  @@  AP  A�  A@  @�  ?�  A  @�  Dv� B�  B,  B�  E�� A�  B  B�  A   A  B  B\  A0  AP  @�  @   @   @   B�  A�  B4  B�  @�  @�  A�  @   A�  AP  ?�  @�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       115L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       s=�k���ӱ@���<�	��9@����@����G!A.�¥R?H[�B�jØ/7�� AH� ��I�3B��Bk��%F�B����WA��N��"�B��6�(��¾���pwAg���� A���M���B��?�\�ǥ�A�I�C.wC���>��»9(BVe�B�9�6��A��0�@�A8X�Bᐆֿ��g@���C��A�.bsa��_���B ��r��¹�Z��M@?�A������5�AhT@�R+�BB�f?��~�!��B �c������o���LA��B���@\�@��nB��/A�;U��8�J���mPGA���³QFB2�H½�g�D�¼eNAܟx�[pA:�:�\d��~%A?��A��9B�/TA�$�	���dA\O�d��BO�WB�.l��WjA�!3�����+م@�D�A�l~�9р�Ҽ`A3�Z@
[����L       
categories[$l#L       *                               	   
                   	   
                  	                                                  
         L       categories_nodes[$l#L                	               !   %   (   .   1   4L       categories_segments[$L#L                                                                                                   L       categories_sizes[$L#L                                                                                                  L       default_left[$U#L       s                                                                                                  L       idi]L       left_children[$l#L       s               	                                    !   #   %   '   )   +   -   /   1   3   5   7����   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c   e   g   i   k��������   m   o����   q������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       sGI}�H4ImHe0>H![5I/�tH�l�H��2HI*H��)I	�H���HH�oI+rlH+� H|UHϝ�I:��HwO'H�`I4HBIqH���I�4H���H��SI7i-H�v!F|    G/^nG�qNH���IJ�GIq8InH�H��mH�֬H�#CH�}�I��H��IR�H���H�3�H��G��H�˔H�,ZH�LH֋HH`�IIyaH�'H��6        F��F���    E�)�                                                                                                                                                                                                                        L       parents[$l#L       s���                                                           	   	   
   
                                                                                                                                   !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   9   9   :   :   <   <L       right_children[$l#L       s               
                                     "   $   &   (   *   ,   .   0   2   4   6   8����   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d   f   h   j   l��������   n   p����   r������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       s>�?}>�S�A         A   >$�/@�  >���   >�o>���?��=� �A�  ?>5?>F��D�@ A  >�  ?L�D@@  >�+>��;>ڟ�         �pw   AP  ??}?A�7   D�@ D�  D��    A0  >��   >�bN@�ƨBD  Bj��>I�^   >�1'@�     @�  >�ȴ   B!  ?Hr���_���A0  BH��¹�ZBG�@?�A������5�AhT@�R+�BB�f?��~�!��B �c������o���LA��B���@\�@��nB��/A�;U��8�J���mPGA���³QFB2�H½�g�D�¼eNAܟx�[pA:�:�\d��~%A?��A��9B�/TA�$�	���dA\O�d��BO�WB�.l��WjA�!3�����+م@�D�A�l~�9р�Ҽ`A3�Z@
[����L       split_indices[$l#L       s                                                  
               
                                     
   
                            
            	                                                                                                                                                                                                                                                                         L       
split_type[$U#L       s                                                                                                      L       sum_hessian[$d#L       sE�8 E�� D�� E�� C�� D�� B   EE  D�� C_  C  D�  C�� @�  A�  E  D@� D�` B�  B�  B�  A�  B�  C�  D�  C	  C&  @@  @   A�  @�  D�� D$@ D  Cb  D#� D?  B�  AP  BL  B�  B�  B  A�  @�  A�  B�  C�� B  B�  D�@ Bx  B�  B�  BT  ?�  @   A�  @�  @   @�  D�� Cy  Ap  D � B�  C� BD  C1  D@ A�  B�  D-� A�  B�  @�  A   A�  A�  A�  B   B  A�  B  @   A�  ?�  @�  @@  A0  A`  A  B�  C(  C=  B  @   A�  BH  D�� B�  B@  A`  B@  A�  B  B�  B   A�  A  @�  @�  ?�  @   @   L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       115L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       ]=A��$��p�B)���'G�2��"'zB�� @f��!2jA�����cO�@������1C��� R��2Aш�Af�9��Aa���
.4�`��B�s�i�A�Q�@}���@�k%��x�C1Bấ��KB2F���B�v�¦ r���u�A�¥ɳ�B���A����A�.�B� �X��@gF�Au	�s~�A�H����A�e@�b��Bf3*���@���B���d��-�3���gBA20DB�ƗB_��uٰA�3��`�{A��jb�A��'��2B�A%AIA6Ԉ��[�Ah6Bö����E�~@�����A=~��;����m&A�@�.P�T���V@g�#L       
categories[$l#L                                             	   
                                     	   
             L       categories_nodes[$l#L       
                     #   +   2   3L       categories_segments[$L#L       
                                                                       L       categories_sizes[$L#L       
                                          	                            L       default_left[$U#L       ]                                                                                L       idi^L       left_children[$l#L       ]               	                                    !   #   %����   '��������   )   +   -����   /   1   3   5   7   9   ;   =   ?����   A   C��������   E   G   I   K��������   M   O   Q   S   U   W   Y   [��������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       ]G���H�fG� fH>nG��VHZ��GuRCHf�PH<�GNP@E̗�G��Hf�I%�H�f�HV[H[��H9�lH\[N    E�7�        G�G��G'Z*    H�0�I0�H�d�H�8�H ��G��E���F�xF�-O    Hmt0H�2�        F��CG�iBG!f�G���        H��IV�I3�KH�eHD��H��TH�H��                                                                                                                                                        L       parents[$l#L       ]���                                                           	   	   
   
                                                                                                                 !   !   "   "   #   #   %   %   &   &   )   )   *   *   +   +   ,   ,   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6L       right_children[$l#L       ]               
                                     "   $   &����   (��������   *   ,   .����   0   2   4   6   8   :   <   >   @����   B   D��������   F   H   J   L��������   N   P   R   T   V   X   Z   \��������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       ]=P�`?�O�=m�h   >���@�        >)��=y�#BD  >�C�   D�� D�@ =ȴ9>^5?D�  >KƨAf@�  Aa���
.4   >�t�A���i�D�  >��w   >�;d=�wA0  D�� >p��   ��>;dZA�  ���u�B[��A�     >��+A����>��#B�  D��       A@  C  ?�O�A�e@�b��Bf3*���@���B���d��-�3���gBA20DB�ƗB_��uٰA�3��`�{A��jb�A��'��2B�A%AIA6Ԉ��[�Ah6Bö����E�~@�����A=~��;����m&A�@�.P�T���V@g�#L       split_indices[$l#L       ]   	      	                  
                        
                                         
          	                                                                                                                                                                                                                                    L       
split_type[$U#L       ]                                                                                   L       sum_hessian[$d#L       ]E�8 B�  Eٸ B�  A@  B\  E�  B,  Bd  A  @@  BH  @�  D�@ E�p B   A0  @�  BH  ?�  A   @   ?�  B   A�  @�  ?�  D/  D�� E+  E	� @�  A�  @�  @�  @@  @�  B  AP  @�  @�  A   A�  @�  A`  ?�  @@  D"� BD  C�� Dx@ D#� E D�� Da� @�  @   A�  ?�  ?�  @�  @�  @   @   ?�  B  @@  @�  A   @�  @   @�  A�  ?�  @@  ?�  AP  C�  C7  B  AP  Ap  C�  D  CЀ C(  C� D�  C  D�` A@  C�  C΀ L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       93L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       �t��n@{'J��/@T�1�}~oA]8|�����p�>ѕBd��
5?�t�B/�懃��]�A˪�'�CD��A>�@�_����`CY~ �A�pBZm"�A�K�o�uBEa����A��B�B����B8`� ��@�'r12C���F�.���B5�e�-R!�+�xÛ��ẠEC��_AS@DAk���̴=³/�B-²6B�rE����A!K���k�B�}B$'�C9�w�V�i@�����3B��y��]�A�<<>/��;oyA�͵�u�F��u[�!�����qA����>J>���C��Aoj��*�.B����@À9A��Q���B"h�Bc����H�ٻ6Aqn�A����|B0rC"��\�'A�2B?��(vAk5����BNg�#�BzՅ?�����B��GB�-A�+��Y~�A.���fA�'�����1ڵBGá����A|�����cB�^���� ��cl�I��A�w���B
@���x��B}�A*��L       
categories[$l#L       ;                         	                           	   
                   	                                           	   
                                     	   
                      L       categories_nodes[$l#L       
   
            %   ,   /   2   ;   <L       categories_segments[$L#L       
                      
                                   +       8       :L       categories_sizes[$L#L       
              	       
                                                 L       default_left[$U#L                                                                                                                  L       idi_L       left_children[$l#L                      	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c   e   g   i   k   m   o   q   s   u   w   y   {   }����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       G}�H:�XHH�`H}�XH�x�H���I	H��dI!�H���I��H�G�H��LI"��H���H��H�A�H��>I=Y�IH
�HԲIbIcP�H�ѲHJ�H���H��H�~�I�rHҍ�HȋH-cH9��I-
6H@/�H���H��PHHG���I�$�I�5I$�$I�LH5��H��IE��H��H�{H���H_�^H�8HAzH���H�N�I0:H��G��ImuI�9_IGVH[�bI	��H�r                                                                                                                                                                                                                                                                L       parents[$l#L       ���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <   =   =   >   >L       right_children[$l#L                      
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d   f   h   j   l   n   p   r   t   v   x   z   |   ~����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       >��yB8  @�  B(G�D�� =�x�>�A�>�-B�  >"��   >ȴ9>�-@   A�           D�  ?gl�>hr�>��>n��B  >�9X=ȴ9>���A   AP  ?��@�  >V>��?���@�  >� �?e��   @�  ?_�w=�x�A\)>j~�B�     >0 �>�A�   D�� D�`    B[��=�S�>��A@  @�  D�@ A   B�        Bu�R=H�9��]�A�<<>/��;oyA�͵�u�F��u[�!�����qA����>J>���C��Aoj��*�.B����@À9A��Q���B"h�Bc����H�ٻ6Aqn�A����|B0rC"��\�'A�2B?��(vAk5����BNg�#�BzՅ?�����B��GB�-A�+��Y~�A.���fA�'�����1ڵBGá����A|�����cB�^���� ��cl�I��A�w���B
@���x��B}�A*��L       split_indices[$l#L                                           	                                 
            	                  
   
            
                                                   	                                                                                                                                                                                                                                                                                               L       
split_type[$U#L                                                                                                                            L       sum_hessian[$d#L       E�8 E�  E$p D�� E D�  D�� D�  C�� E� C  CO  D�@ D
� D  D*� DW� C�  A0  D�� D�  B�  B  C   B�  B�  D�� Bx  C�  C�  C  B�  D@ C�  D	� C  CP  @�  @�  DY� C� C�� D6� A   B�  A�  A`  B  B�  A�  B|  A`  B�  C�  D4� B@  A`  C� A�  CP  Cz  B�  B�  A`  B�  C(  C؀ C#  C  D� A0  A�  B�  C  Bd  @�  ?�  @�  @   DT� A�  C�� C(  C�  A�  Ap  D2� @�  ?�  B�  A�  A@  A   @�  A   A  A�  A`  B�  @   A`  A   B\  AP  ?�  @@  B�  C�� B�  D� B�  A�  A�  @�  @�  CЀ B@  A�  @   C!  B<  B  CT  BP  AP  A�  B�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       127L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       I=&�A���S�2�n�pB����2�o���B����</5B��'����l�Ba �BT��[�Bh�B����BO,�C1�t@��U�1���Q-@䡦C0�[�4k�	��BKKM@gh BC��k�A�U~�_^gA��C�o~�H�B�
�@��D°� BA����$zB���Al��(�c��AB�l�CA�M@��g@^6��(A���?����f�$�E��A0�B�}��3�A_́�^T�A������AX^���s�A�� B�7��]�
g4���?@"AлTA�������L       
categories[$l#L                                             	   
            L       categories_nodes[$l#L                   ,L       categories_segments[$L#L                                    L       categories_sizes[$L#L                                   L       default_left[$U#L       I                                                                   L       idi`L       left_children[$l#L       I               	               ����   ����         ����         !   #����   %   '   )   +   -   /   1   3   5������������   7   9����   ;   =   ?   A������������   C   E   G��������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       IGT��Hw?Gh�G��G���GڳRG��,FE� G��H��    G�G�    HH�H][,E6�\    G�yE�ҔG�E�H ��    GG�G �F���GM��Gr��B,5 C�(EZdG4�0            G�<�Ga�6    G2ƼF�F�jaGHdj            E�0H���G�>v                                                                                                        L       parents[$l#L       I���                                                           	   	                                                                                                         "   "   #   #   %   %   &   &   '   '   (   (   ,   ,   -   -   .   .L       right_children[$l#L       I               
               ����   ����         ����          "   $����   &   (   *   ,   .   0   2   4   6������������   8   :����   <   >   @   B������������   D   F   H��������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       I<�C�B   <���Ap  D�� @n�D�  D�  A   Bb  ���>!��Ba �>�G�D�` >�(�B��>+B�  >�O�B�  �1�@@  >P�`B`  >�1'D�`          BH��A�U~�_^gA��B2  ?�=qB�
�B!  >���B�  A�  B���Al��(   @j�H<oA�M@��g@^6��(A���?����f�$�E��A0�B�}��3�A_́�^T�A������AX^���s�A�� B�7��]�
g4���?@"AлTA�������L       split_indices[$l#L       I                  
                                	                          	                                                                                                                                                                                       L       
split_type[$U#L       I                                                                     L       sum_hessian[$d#L       IE�8 B\  Eۀ A�  A�  A�  Eژ A   A�  A�  @@  A�  ?�  A�  E�� @�  @   A�  @�  AP  A   @�  A�  A�  @�  @�  E٠ @�  @   @@  Ap  @�  ?�  @�  @�  @�  ?�  A`  A   A  A   @�  @   @@  @@  CĀ E�X @@  ?�  ?�  ?�  @   ?�  A  @�  @   @�  @�  @@  @�  @�  @�  ?�  @@  @�  ?�  A  ?�  @   C�� B8  B   E� L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       73L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       m=�-�@$�M�1��@K���.A0{r�
�?�k�B����r���3�k׫B3������@�@j�����_A�B�K������8�����B�$AY��'ʒA<��B���AsA����B��:4@��?@:rTC	@2�xh-�1S©�_B�4�B���6)ȿ���������հ�@`6��pB;���QR EA�U�CZ�@�jC"?S�z��B����/`B��I�/��E?�vbBU|L?��?��d������UMB�����]B�ý�k���L�-� ��@<�B�BP?7�)BT�JB�ˇ��V�
X�@�agBEc�@�y�raAM�VB:����*�����B%��A���f&_A��B�0��DXyA�L�Bh���
kA��m�
�B�6�@�����]���A�;D��Il�Aͅ�mA����e�`	?��L       
categories[$l#L                          
                               	   
                           L       categories_nodes[$l#L                   "   #L       categories_segments[$L#L                             
              L       categories_sizes[$L#L                            
              L       default_left[$U#L       m                                                                                                  L       idiaL       left_children[$l#L       m               	                                    !   #   %   '   )   +����   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K����������������   M����   O   Q   S   U����   W   Y   [   ]   _   a   c   e   g   i   k������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       mGD�$H7eH���H`>�H��H�"WH֓0H�GQH�dGI8�F�H�N:I&f`H��H�дH�zGH��HT4�H��.C�?(F�PF�Z    H�k�H�-�I�SIP/�H��@Ib�cH��~H`�(HY$MIZ�H��%H�+�H��G�>�I(PHI�6                FG    I2�H�/�H��dH��n    H���I�(H�;H�
H�Z H*�I[��H�_I3^?H�Q�H[�<                                                                                                                                                                                                L       parents[$l#L       m���                                                           	   	   
   
                                                                                                                                   !   !   "   "   #   #   $   $   %   %   &   &   +   +   -   -   .   .   /   /   0   0   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <L       right_children[$l#L       m               
                                     "   $   &   (   *   ,����   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L����������������   N����   P   R   T   V����   X   Z   \   ^   `   b   d   f   h   j   l������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       m@aG�?f$�D�  ?ƨ?�m@�  D�  >�x�D�  B'
=B�  D�` D�` >>v�>�b?�^5?oA0        @�  @,�B�$@   @�HD�` >��F@@  @�  @�     ?��B0  ?M�      ?�(�B33=�^5����������հ�?�o�p>��@�>)��>�bCZ�?I�?���?2-?)�^=��?�#B�  >%�TB�33?'l�@qG�?��d������UMB�����]B�ý�k���L�-� ��@<�B�BP?7�)BT�JB�ˇ��V�
X�@�agBEc�@�y�raAM�VB:����*�����B%��A���f&_A��B�0��DXyA�L�Bh���
kA��m�
�B�6�@�����]���A�;D��Il�Aͅ�mA����e�`	?��L       split_indices[$l#L       m                                                   	                                                       	                 	                   
       
      
                   	            
      	                                                                                                                                                                                                   L       
split_type[$U#L       m                                                                                                        L       sum_hessian[$d#L       mE�8 Ej� EO� Ei A�  Dx@ E� E^� C$  AP  A`  D-@ C�  B�  E
� ES` C7  B  B�  @@  A   AP  ?�  D   C5  CK  B�  B$  B�  Dz@ D�� ER@ A�  C  B  B  @�  B�  B4  ?�  @   @�  @�  A0  @   C"  C�  B�  B|  ?�  CJ  B�  A�  A`  A�  A@  B`  DG� CJ  B�  D�� E0� D� @�  A@  C  @�  A�  A�  A�  @�  @@  @   A�  BL  @   B,  @�  @�  B  C   Ct  B�  @�  B�  B0  A�  B   C"  B  B  AP  A   A0  @@  A  A�  @�  @�  B  A�  B�  D6� C5  A�  BH  B,  B�  D�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       109L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       a=�x6����@�����>��n�C&s�@,?13���0B�s��o�DEH�B�$�@MR��D2@�
��A7���2��A�����CBy���A��oC��PA�� �"C��A ���ՆA� '��\ �X^!A����ft���5�ĸB�y���m/A�w���3Cv�*_��|]~C5 0�6bi�z�U�Cup�vs@�qB�8�怚������<�@uB��4�ҙ-��GbA��>�a��9��������n�A�m�@��B��jA� �$f��͋�@;4Aߊ�B��BA[��������ŉ�B��'�l#4��n?�Kg?yT� ]gB���C�M����A�A@)���o BE���������@�2@ɻHڋL       
categories[$l#L       &                                                                            	   
                               
         L       categories_nodes[$l#L       	            $   &   +   /   1   4L       categories_segments[$L#L       	                                           	                     L       categories_sizes[$L#L       	                                                               L       default_left[$U#L       a                                                                                     L       idibL       left_children[$l#L       a               	                                    !   #   %   '   )   +   -��������   /   1   3   5��������   7   9   ;   =   ?   A   C   E����   G����   I   K   M   O   Q   S����   U   W   Y   [   ]   _������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       aGTńH�y�I.N�G�RbI!y
I�҄Hh~H1�H!~�H[��H��I��H���HF��G�@�H�H��HYo H"-Gc��H�VH�ȜH��i        G<�H���HN�H�\�        H,�I�nH���I��HT�.H�xH6�H�1    Fy�    GZ�`H6�XH�� G�<,H;2*D2��    HY�tG:��HRVdH�=H�mbI/_                                                                                                                                                                        L       parents[$l#L       a���                                                           	   	   
   
                                                                                                                 !   !   "   "   #   #   $   $   %   %   &   &   (   (   *   *   +   +   ,   ,   -   -   .   .   /   /   1   1   2   2   3   3   4   4   5   5   6   6L       right_children[$l#L       a               
                                     "   $   &   (   *   ,   .��������   0   2   4   6��������   8   :   <   >   @   B   D   F����   H����   J   L   N   P   R   T����   V   X   Z   \   ^   `������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       a>�>�V>�Q�?1'@   ?�
@�  >\@�  ?CS�A  B̊==�h@�     >���?Rn�@�  ?�{   >$�/Bb  D�� C��PA��    >�5?A0  A�  A� 'D�` >VD�  Ap  @@     D��    A�D�` ��3B     >�=q@��R@�     �   >ؓuB�=q   @s33?Y���<�@uB��4�ҙ-��GbA��>�a��9��������n�A�m�@��B��jA� �$f��͋�@;4Aߊ�B��BA[��������ŉ�B��'�l#4��n?�Kg?yT� ]gB���C�M����A�A@)���o BE���������@�2@ɻHڋL       split_indices[$l#L       a   	   	   	                     
                     
                                                     
                                        
                                                                                                                                                                                                          L       
split_type[$U#L       a                                                                                        L       sum_hessian[$d#L       aE�8 E� D�� E�x B�  A�  Dŀ E�� Cs  A�  B�  @   A�  D�� @�  E� D�@ C  B�  A   A   BH  A`  ?�  ?�  @�  A�  D�� Cq  ?�  @�  E|� Bh  DU� CD  B�  A�  AP  B�  @   @�  @   A   A�  A�  A   @�  @   @   A0  A  D�  B  CJ  B  EO� D4  @�  BT  CJ  D#  C(  A�  B�  A�  @�  AP  A   @�  A�  B|  @�  ?�  @@  @�  A@  A�  @�  A`  @�  @   @@  @@  ?�  ?�  A  @   @�  @�  D�� B�  A�  A`  B�  C  A�  A�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       97L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       i=�h|��A�j���%`�BfX�.l��Қ�?ө[B8�à*vA��OC	n��A�bo�5�>��C�?�#�Bz[gA&�w��@�B�AAg�VCg*�CA����UpA�@Ç�xCN�� ���eD&B�>RA.��C��9A��=<�9B"y�B� ������X}���Z�5�B�2B��NA��Bv(�C��NB(���)���0��Bk �����s�C��	��q ôE��@2_��C�����B�-G��N��)��A��n5AB5�C�9�ֳ\BCjp>�X-����A��;��^�@4B��]��@�4��.� �.�	� +A��B�"@���B=�4?ק4C�B-i�A�[T�9��@��� �����r���`��A�B�PA�CB�����i�-O��ٜA����iL       
categories[$l#L                                         	   
                 L       categories_nodes[$l#L                3   9L       categories_segments[$L#L                                    L       categories_sizes[$L#L                                   L       default_left[$U#L       i                                                                                                  L       idicL       left_children[$l#L       i               	                                    !   #   %����   '   )����   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O����   Q   S��������   U   W   Y����   [����   ]   _   a   c   e   g����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       iG��G�7lH�=�G�+�I0�Hw�H���HW#H�ەG��I~��H^��He�H���I>X�H�m�I	�\IH�>HN�$    G)>ZH��    HX,�G,��H� ~G�6G)VH�A�H��VH�
�H�xIB��I��I!qFH��H��iH �OI'��F�|Fo��F�o�    H�K�H�3�        GdTqH�(F�    E��    I��G��0G‰H|�aH|G�q	                                                                                                                                                                                        L       parents[$l#L       i���                                                           	   	   
   
                                                                                                                             !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   +   +   ,   ,   /   /   0   0   1   1   3   3   5   5   6   6   7   7   8   8   9   9   :   :L       right_children[$l#L       i               
                                     "   $   &����   (   *����   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P����   R   T��������   V   X   Z����   \����   ^   `   b   d   f   h����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       iB�  Bճ3D�� >�"�?vE�D�� @)��>��>�(�=�j@BM�B�  @�  >O�>�|�>��\>bN=�Q�B�ǮBz[g=�%   B�A=�9X   >�
=@�  ?.{>ٙ�@�{>��>�-@�  BT  D�� =0 �>��TB��{@��@�  ?$Z@   ���Z>�I�=�Q�B��NA��>��B�  @�  �)��   Bk =�S�@@  >��=�-   ?�@2_��C�����B�-G��N��)��A��n5AB5�C�9�ֳ\BCjp>�X-����A��;��^�@4B��]��@�4��.� �.�	� +A��B�"@���B=�4?ק4C�B-i�A�[T�9��@��� �����r���`��A�B�PA�CB�����i�-O��ٜA����iL       split_indices[$l#L       i            
            
   
   
            	      
                                                                                        
                                  
      	                                                                                                                                                                                                 L       
split_type[$U#L       i                                                                                                     L       sum_hessian[$d#L       iE�8 E�� C�  E�@ A�  CM  Bl  D�` E�� A�  @�  C6  A�  A�  B  D�  C�� A�  E�� @   A`  @�  ?�  C2  @�  A�  @�  A  A`  A�  A�  D�� A�  C  C"  @�  A�  E�� C  @@  A0  @�  ?�  B4  C  @   @   A   @�  @�  @   @�  @   @�  A   A@  A   @�  A@  DL@ C�  A�  A0  B�  B�  B�  B�  ?�  @�  A   @�  E�  C�  B�  A�  ?�  @   @�  @�  ?�  @�  A�  A�  @@  C  @@  @�  @@  @@  @@  @   @@  @�  @   @   @�  @@  A   @�  @   @�  ?�  @@  @�  @�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       105L       size_leaf_vectorSL       1}}}L       nameSL       gbtree}L       learner_model_param{L       
base_scoreSL       3.7122964E3L       boost_from_averageSL       1L       	num_classSL       0L       num_featureSL       24L       
num_targetSL       1}L       	objective{L       nameSL       reg:squarederrorL       reg_loss_param{L       scale_pos_weightSL       1}}}L       version[#L       ii i}}�
       ���R�sbub.