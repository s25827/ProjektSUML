��/      �xgboost.sklearn��XGBRegressor���)��}�(�n_estimators�N�	objective��reg:squarederror��	max_depth�N�
max_leaves�N�max_bin�N�grow_policy�N�learning_rate�N�	verbosity�N�booster�N�tree_method�N�gamma�N�min_child_weight�N�max_delta_step�N�	subsample�N�sampling_method�N�colsample_bytree�N�colsample_bylevel�N�colsample_bynode�N�	reg_alpha�N�
reg_lambda�N�scale_pos_weight�N�
base_score�N�missing�G�      �num_parallel_tree�N�random_state�N�n_jobs�N�monotone_constraints�N�interaction_constraints�N�importance_type�N�device�N�validate_parameters�N�enable_categorical���feature_types�N�feature_weights�N�max_cat_to_onehot�N�max_cat_threshold�N�multi_strategy�N�eval_metric�N�early_stopping_rounds�N�	callbacks�N�_Booster��xgboost.core��Booster���)��}��handle��builtins��	bytearray���B�n {L       Config{L       learner{L       generic_param{L       deviceSL       cpuL       fail_on_invalid_gpu_idSL       0L       n_jobsSL       0L       nthreadSL       0L       random_stateSL       0L       seedSL       0L       seed_per_iterationSL       0L       validate_parametersSL       1}L       gradient_booster{L       gbtree_model_param{L       num_parallel_treeSL       1L       	num_treesSL       100}L       gbtree_train_param{L       process_typeSL       defaultL       tree_methodSL       autoL       updaterSL       grow_quantile_histmakerL       updater_seqSL       grow_quantile_histmaker}L       nameSL       gbtreeL       specified_updaterFL       tree_train_param{L       alphaSL       0L       	cache_optSL       1L       colsample_bylevelSL       1L       colsample_bynodeSL       1L       colsample_bytreeSL       1L       etaSL       0.300000012L       gammaSL       0L       grow_policySL       	depthwiseL       interaction_constraintsSL        L       lambdaSL       1L       learning_rateSL       0.300000012L       max_binSL       256L       max_cat_thresholdSL       64L       max_cat_to_onehotSL       4L       max_delta_stepSL       0L       	max_depthSL       6L       
max_leavesSL       0L       min_child_weightSL       1L       min_split_lossSL       0L       monotone_constraintsSL       ()L       refresh_leafSL       1L       	reg_alphaSL       0L       
reg_lambdaSL       1L       sampling_methodSL       uniformL       sketch_ratioSL       2L       sparse_thresholdSL       0.20000000000000001L       	subsampleSL       1}L       updater[#L       {L       hist_train_param{L       debug_synchronizeSL       0L       extmem_single_pageSL       0L       max_cached_hist_nodeSL       18446744073709551615}L       nameSL       grow_quantile_histmaker}}L       learner_model_param{L       
base_scoreSL       8.2300875E5L       boost_from_averageSL       1L       	num_classSL       0L       num_featureSL       24L       
num_targetSL       1}L       learner_train_param{L       boosterSL       gbtreeL       disable_default_eval_metricSL       0L       multi_strategySL       one_output_per_treeL       	objectiveSL       reg:squarederror}L       metrics[#L       {L       nameSL       rmse}L       	objective{L       nameSL       reg:squarederrorL       reg_loss_param{L       scale_pos_weightSL       1}}}L       version[#L       ii i}L       Model{L       learner{L       
attributes{}L       feature_names[#L       SL       citySL       typeSL       squareMetersSL       roomsSL       floorSL       
floorCountSL       	buildYearSL       centreDistanceSL       poiCountSL       schoolDistanceSL       clinicDistanceSL       postOfficeDistanceSL       kindergartenDistanceSL       restaurantDistanceSL       collegeDistanceSL       pharmacyDistanceSL       	ownershipSL       buildingMaterialSL       	conditionSL       hasParkingSpaceSL       
hasBalconySL       hasElevatorSL       hasSecuritySL       hasStorageRoomL       feature_types[#L       SL       cSL       cSL       floatSL       floatSL       floatSL       floatSL       floatSL       floatSL       floatSL       floatSL       floatSL       floatSL       floatSL       floatSL       floatSL       floatSL       cSL       cSL       cSL       cSL       cSL       cSL       cSL       cL       gradient_booster{L       model{L       gbtree_model_param{L       num_parallel_treeSL       1L       	num_treesSL       100}L       iteration_indptr[#L       ei iiiiiiiii	i
iiiiiiiiiiiiiiiiiiiiii i!i"i#i$i%i&i'i(i)i*i+i,i-i.i/i0i1i2i3i4i5i6i7i8i9i:i;i<i=i>i?i@iAiBiCiDiEiFiGiHiIiJiKiLiMiNiOiPiQiRiSiTiUiViWiXiYiZi[i\i]i^i_i`iaibicidL       	tree_info[#L       di i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i i L       trees[#L       d{L       base_weights[$d#L       �O�F���=Ic�EF�>ȯ�MIQŗF�q�Ƕ�H2b��к��y�I�I��HR��Ƕ���=����H�c�Gդ�Ȥ����,Ȕ���ج�I.��H�pWI���In��G�>fH�����G#Ԕ�ό�j@�F'u��˷Hʚ�GD��H2�����ȳX{ȃo)��s]Ȭ=��kkTȫ�
ƬIq��IBIT��I	BDHo(]I���I���I���I�&G=�H��H���H=��!�C��G❒�[?(ƴ�P�T7��OǞ�G2����9y�FC�F	HG���H�Gf	wƟ��F���G��@ƄEG �������<���^�Ǆ�Q�C �_��TgǫK��L&tǜ�Җ��9�L�nE���n*����H#��Hj�H�\#H8�H;�|G��6G�vIG&��H��#H�J�H�x�H�Q
H�H�H�?H
��Hx��F�U��+hG�tGdYG�X�H
�G�$�G
�~�v]�.�F�d��f�G��hF���ś���#L       
categories[$l#L       �                      	   
                            	   
                                        
                        
                                               	   
                                     	   
                        
                      
                               	   
                                            	   
                         
                                                      	   
                                     	   
                     
                
L       categories_nodes[$l#L                      	                                       "   $   +   ,   /   0   2   <   =   >L       categories_segments[$L#L                      
              !       "       '       (       ,       /       :       G       L       S       T       a       b       p       u       v       w       {       |       }       �       �       �       �L       categories_sizes[$L#L              
                                                                                                                                                                                      L       default_left[$U#L                                                                                                          L       idi L       left_children[$l#L                      	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c   e   g   i   k   m   o   q   s   u   w   y   {   }����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       XlV�W�%W�[bW"2UݔpV�ȰU�ԛV=�VD�U��U1O�U��PU�6�TD�Tt�T���U��BU���U���S�T@TE�TWM�S���U� T`2T��UC1�S��ZS~s�S���S/�T;�T��U\�T��T�Q TZ�U6��T���S;�SN S�G S	� SHc S`J�R�fS�8T��T��@S0j@T��Ta@Tr�U {�T/0R��;R�~�R��`R�c�S R��R���Q��                                                                                                                                                                                                                                                                L       parents[$l#L       ���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <   =   =   >   >L       right_children[$l#L                      
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d   f   h   j   l   n   p   r   t   v   x   z   |   ~����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       B�ff      B\  BT��B�(�   B�R      D�� ?�S�   B�  D��             D�` D�        B�     A�           B�     @\��@�\@G
=   B�     B�  B�\B(  B\)B#
=B.��      Bi��Bt        @?;d   B�  B�  @p�B�  A0  ?$��D�  >�C�B�           ƴ�P�T7��OǞ�G2����9y�FC�F	HG���H�Gf	wƟ��F���G��@ƄEG �������<���^�Ǆ�Q�C �_��TgǫK��L&tǜ�Җ��9�L�nE���n*����H#��Hj�H�\#H8�H;�|G��6G�vIG&��H��#H�J�H�x�H�Q
H�H�H�?H
��Hx��F�U��+hG�tGdYG�X�H
�G�$�G
�~�v]�.�F�d��f�G��hF���ś���#L       split_indices[$l#L                                               
                                                                                                                             
                                                                                                                                                                                                                                                                                                          L       
split_type[$U#L                                                                                                           L       sum_hessian[$d#L       F�` Fc� E$ F P E�� D�  D^  E�X E`� E#� DӠ D�  D2  C�� D� E� E�h D�� E� DW� D�� D�  Cڀ DO  CE  C�� C�� C  CR  Cր B�  D�  D�� E4 D�� Da� CW  D�` Dp@ D  C�� D�� C`  D� D4� B�  C�  D� C�� BT  C  C  CQ  C�� B�  B�  A�  C	  B�  C�� B�  Bh  B0  C�  D@� CĀ DG  D� E� D�  Cd  C�  C�  B�  B�  Da� D  D(� C�� CL  C�  B�  C3  D!  D^� B�  B�  C  C�� D-� A�  A�  B�  B�  C7  C�� C  C�� B  B  Ap  BP  B�  B�  B�  B,  C&  B�  C3  BX  B(  B�  A0  A�  A@  B�  A�  B  B  C  C-  B  B�  A�  B(  A�  A�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       127L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       C<��Ǘ�|H�Y��CEG�yuItWFb.ǮC�G��Ȑ���+BKH�eeI]fOH��Ǎ�\���[N9HS.ņ��dyȠ��H��i�7I	q�H�DdIy��I+g�G�-VHL��Ǻ^TF欇��ɛ�V0��q�q�о H��<G��ǝn$G֗��w���)H?ȦO�k������h�tƛ��ӟ[H�rI1�HM�`H��I�TjIS@0IX�IGF{�HE��H�ZEH&�4��`-C=�G�|��;�Lk8�+i�;4�ǌl��*9�F�{��+ �Ƒ{2Gf�G� F5�hGI�G���ڡ�G˓[F��ǭaǉ!�ǉ��� _��s�Ƕu�Ǹ��t<k�����O�yǚ���Z%d�S,VF��t���Aǃ�QH,rG��HiK�G���G�|2G&��HKVLG��H���H���HW��H��HZ��G�s>H� �H7��}F���G�E�ſ1�G2�JG�=^F�_G����}�&A/��QF��G�C���ƌȤFI��L       
categories[$l#L       �                      	   
                            	   
                                        
                                  	   
                        
                        
                
                                   	   
                                          	   
                                    
                                  	   
                                        	   
                                            	   
                         
       L       categories_nodes[$l#L                      	                           !   +   -   .   0   1   5   7   8   ;   =L       categories_segments[$L#L                      
              !       .       3       6       ;       @       A       O       P       Q       ]       ^       b       c       e       f       t       �       �       �       �L       categories_sizes[$L#L              
                                                                                                                                                                 L       default_left[$U#L                                                                                                     L       idiL       left_children[$l#L                      	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c   e   g   i   k   m   o   q   s   u   w   y   {   }����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       W�cW+��W>��V��}UJ�Vz�`U%�^U A�U���T�Z�T��`U���U� S�{pS��TpT�@"U�TUh�hSyX�S�� Sɡ�Sn|U@U��T{� T/� S���S;<�S��(R�S��R�^@T�`�T��U&�UW�T�T�1�R� S��S�� R�`RƟ`SCQ R�jR���T��T���TάT+��S�� Te�S�1S֡@R��vR��R8��SD��R�,PR�<R2nQ��L                                                                                                                                                                                                                                                                L       parents[$l#L       ���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <   =   =   >   >L       right_children[$l#L                      
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d   f   h   j   l   n   p   r   t   v   x   z   |   ~����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       B�        BH  B[z�B�     B        D�� ?VE�>k�B�  D�     ?BM�@~{D�  D�` D�`       B�           D��    B�     ?��?��R   D�� Bq33Btp�?�R?���B(  B&ffB-��B\)   B���      @qG�      >+@��D�@    ?�+      D�� B�     ?+ƨ   @��R�Lk8�+i�;4�ǌl��*9�F�{��+ �Ƒ{2Gf�G� F5�hGI�G���ڡ�G˓[F��ǭaǉ!�ǉ��� _��s�Ƕu�Ǹ��t<k�����O�yǚ���Z%d�S,VF��t���Aǃ�QH,rG��HiK�G���G�|2G&��HKVLG��H���H���HW��H��HZ��G�s>H� �H7��}F���G�E�ſ1�G2�JG�=^F�_G����}�&A/��QF��G�C���ƌȤFI��L       split_indices[$l#L                                                
                
                                                                                                                                                                                                                                                                                                                                                                                                                    L       
split_type[$U#L                                                                                                              L       sum_hessian[$d#L       F�` F_p E5@ F` E�  D�� D{@ E� E�� E-� D�` D�� C�  Cɀ D� D�� EW� E:� D�  Dg� D�` D�` C�  Db� C�� C�  C0  CA  CR  C�  B�  D�� C� D� D�� DT� E� D�` D7� D-@ Ci  D�@ Ci  C�� D%� C#  C  D� C�  C�� C  C/  C  B�  B�  C  Bh  B\  C  C�� B�  Bt  BD  CS  D�� B�  C�� D�@ C�� DL� D3  C�� C�  D�  DT� B�  D�  B�  D� CV  C� B�  C  DM@ DG@ B�  C#  C  C�� C�  C\  B�  B  B�  A�  C�  C�  Cf  Bh  C  CX  BT  B�  B�  Bp  B�  B@  A�  B4  B�  A�  B�  B�  BD  A  A  B8  B�  B�  B�  C�  B�  A�  B  A�  B  A`  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       127L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       C��Ǉ��HUVq�a���_�H����qBǐ�^G07o�рh�J��Hpm�I�YG�˟�A�6�6��ǹlnH�E��Y�f�ǆPD�[�F��MH:��H��Ie"H�g5G��,H;��ǟJ�EI�Lǩ��F[ɥ��"ǔۭH3��Gp.�H	�ş,�,�-��Iǻ��FS[��p�\�@���CX���:eHpGG�8'H�V IuI56�I ��H��(I|�Fӊ H��H�vH�� �ߒe��G]1��'��$���6����=F�܍�GO_��;EВ����KF�?�G}J�F����P��Gn�jF�ICF;��i���Z�P�#r8F+�q�%6ŷ�/��Z��?�G��qǣ�ǈy��[A�ǓLǈ���OY>�����0AG�FLF�ظF�>G���G�X�F���H@�G�n	F�6�H\ jHd�H��G��EGMG�j�H<��G��mE���G�	�F�@F�5HG����{:�G�I�ƫȆ�(?`E�_�Ƣ��E�&+GH';Řy����'L       
categories[$l#L       e                         	   
                               	   
                            
                                  	   
                                          
                                   	   
                     
                                	   
                         
               
            
L       categories_nodes[$l#L                                     $   %   &   ,   .   1   5   ;   <   >L       categories_segments[$L#L                                           ,       -       .       /       0       6       7       E       G       I       J       W       X       ]       bL       categories_sizes[$L#L                                                                                                                                            L       default_left[$U#L                                                                                                          L       idiL       left_children[$l#L                      	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c   e   g   i   k   m   o   q   s   u   w   y   {   }����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       Wn6�V�'�V�{RU�)�UO��VMN(T�5TS��U���T��T1c`U_,�U#6pS�v S�a<S�=�S��@T@�hT�_S�׀TI+@S�A@S5��T�T�T�] T�� T�a�Sx��R���SstSt��R�H,S?wRP?�S�HT� S���Sv �T���R�� S��SK�0S��R� R�S Q׽�R���T�0 T9�TO
`S'��S�� T�/�TNP�Sx4@R�j�S�RйR
�PR���SohS!��Rp<&                                                                                                                                                                                                                                                                L       parents[$l#L       ���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <   =   =   >   >L       right_children[$l#L                      
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d   f   h   j   l   n   p   r   t   v   x   z   |   ~����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       B�        B.��   B��         B@��D�  A�  >k�B�  D�  BffB��>�J@z�D�� D�� B@  B-��   D�     B�  D�� D�� B��{   @�  B<  A�  @	��BC��         B:ff?c�
?��A�  B��   B\)   @�jD�@    >ۥ�=�>�   >�V>�Q�@VffB�  =��
      B�     �$���6����=F�܍�GO_��;EВ����KF�?�G}J�F����P��Gn�jF�ICF;��i���Z�P�#r8F+�q�%6ŷ�/��Z��?�G��qǣ�ǈy��[A�ǓLǈ���OY>�����0AG�FLF�ظF�>G���G�X�F���H@�G�n	F�6�H\ jHd�H��G��EGMG�j�H<��G��mE���G�	�F�@F�5HG����{:�G�I�ƫȆ�(?`E�_�Ƣ��E�&+GH';Řy����'L       split_indices[$l#L                                                                                                                                                               
          	      	                                                                                                                                                                                                                                                                                                 L       
split_type[$U#L                                                                                                                   L       sum_hessian[$d#L       F�` FK� E�@ E� E�� E$� D�� E.� E�X E+� E7P D�` D[� Cɀ D�` D/  E� D�� ES� D�` D�@ EP D(  D�@ C�� D	� C�� C�� B�  D0@ C�  C2  D� D� D�  DX� C�  C�� E@� DT  C�� D�` C�� D�� Dt@ CL  C�  DO@ C� C�  B�  C�  C|  Cb  B�  C5  B�  B�  A�  Cˀ C�  CE  Ce  B�  B�  C΀ B�  C\  C�� C:  D�� Cb  D @ C[  B�  C  C&  D�@ D�  D&� C5  A�  C�  C  D� C�� A�  C�  De� DN@ C  B�  B�  Ce  Co  D$� C*  C�� B�  C�  B0  B�  A�  @�  C�  Bd  CC  B�  B�  AP  B�  @�  C/  B0  BP  B@  B<  ?�  A�  C*  Cm  B�  CD  C  B$  C  B�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       127L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       }C�K���H]BDF�K���"PH���G���ƌ=DG�&��r]�)�zH���HG`+H�"���G&���H�G&��ǰ�!��<ǑGvF�CH�H��H�AH�
{G�h�Ho4�ƛ�G�n��t��G��Ǉ��\�H;��Gl�F��G���D{�<O������r�ƲZ&��I�G��;���I:nH��'HT�IGҏ�H��OH�ّHO��G"�HeɑH���H��GȞ��+H6�rG��>�%�#FH[F��~G]���V>���{���v�F�^*G���G�F]ՅG���G)/�D�:G��E���ʾƦ5�ʮ�����8&��q o�<���肞Fup�6���1F!�:G�*`Ff�$��0\��ւH\;HK.�G��Hc2G�1�F�-�G�T�H0��G���F��6G���G�/G���FqS�F��_�K�F]=GG��$G���G(F��G��Ƒ)iF�kq������E�Gm҂F��nŵ�
L       
categories[$l#L                                	   
                                     	   
                                     	   
                                     
                                    
                                  
                                        	   
                            
                                  	   
                
          
                            	   
                L       categories_nodes[$l#L                            	                        #   )   ,   .   7   9   <L       categories_segments[$L#L                                           &       '       (       0       1       2       <       H       V       ]       j       k       m       n       p       q       ~L       categories_sizes[$L#L                                                                             
                                                                             L       default_left[$U#L       }                                                                                                    L       idiL       left_children[$l#L       }               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c   e   g   i   k����   m   o   q   s   u   w   y   {��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       }V�	�V8ӽV;�^U�BkU��U6d�T�{�T�z�T�+\T�QPT�9(T�� To֜Tn��S�TV-TD;�Tf��S��
S�pS;�S�FTf%T�o`T��S��8S���S�f�T'T�R���Q���S'b�S���S��hT0?TS2=2S��@Te0@S�SuP�R�Rt R���S!p TV�R�xS���T_�`SF\�S� S��S�lS2X    SC�hR���Sѐ�S��`R�RYR�$�P�E Q���                                                                                                                                                                                                                                                        L       parents[$l#L       }���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   7   7   8   8   9   9   :   :   ;   ;   <   <   =   =   >   >L       right_children[$l#L       }               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d   f   h   j   l����   n   p   r   t   v   x   z   |��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       }B��      Bg��Bh                 D�  @��B�ff      B(��B)�@n�D�� D�� D�           B�  D�  B  B�  >_;d      @�  B8  @�=qA�     ?�9X@�\?|�@@  @���   B�R?�z�   ?��
   >�bNB  ?�/?���@~{?q�>�VHO��   >6E�   B���>"��   >�Q�?�h�%�#FH[F��~G]���V>���{���v�F�^*G���G�F]ՅG���G)/�D�:G��E���ʾƦ5�ʮ�����8&��q o�<���肞Fup�6���1F!�:G�*`Ff�$��0\��ւH\;HK.�G��Hc2G�1�F�-�G�T�H0��G���F��6G���G�/G���FqS�F��_�K�F]=GG��$G���G(F��G��Ƒ)iF�kq������E�Gm҂F��nŵ�
L       split_indices[$l#L       }                                                                                                                              
                                            
              	                                                                                                                                                                                                                                                                           L       
split_type[$U#L       }                                                                                                        L       sum_hessian[$d#L       }F�` Fh� E F� E̠ D�` D�� E�0 EP E�  E@ DU� C�� D
� D  D�� E�� D�� D�  D�� E� D�� D  D� C�  C�  BD  C�� C�� C�  B8  D� DQ� D�@ E$� Dt@ C�� DJ� C~  D�@ D	  E� CȀ C�  Dw  C�� C�� C�� C[  CK  B�  CH  B�  B  A`  Cy  B8  B�  C  C  C�  A0  B  C�  C  D1  C  D{� Dd� E` C�� D� C�  C�� A�  B|  D;  B�  C  D�� C�� C�� C�� D�� C�� B�  C�  BH  C�  Dm� B  BX  C�� C  A�  C�  B�  C  B�  C'  B  A�  Bp  BX  C  B,  B  A�  @�  C*  B�  A0  B  B�  A�  B�  B�  A�  B�  C�� Bl  ?�  A   A�  A  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       125L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       C������G�4�F�d��f�HY�F��1�J�kG�F�ǟ���t�,H#��H���ƀ�G�F)���8$�HIF����s����|��,��F��%H|��G�a:H�:Hs��F����0{6H0{MG���(��G��Ǉ��JzaG�y�H��G��9zG�*�ǆt"F'���.��
hEǔ�\ƪY G����&	H��IH({�G'��HiH�A�I��H�O�H?�	CQ�RG�� ���n�H���G�bG�����Ƥ��D�L����G(qƒf���YZ�1�	F�"GL�DF��G�ݭE��|D��=ƥi�F�4���|L���tJ�ſ�F�j�����&j�(u��B��S�C�ݓ��T2;Ǝ �G�rF	��Ƌ۳En1�G��G{�����uG_aF�wmƃ~�G\��Ž�G"Y'G���H(u�G5��H!F���H
�dGE�c�&�gG�OF�\�G��\�3~�F����/���{���^mG�G5����i9F�9O�?V\��i�F� cL       
categories[$l#L       n                               	   
                                     	   
                            
                        
                               	   
                                      	   
                                           	   
                                            
                                    	                L       categories_nodes[$l#L                	                           !   %   +   2   9L       categories_segments[$L#L                                    "       #       +       8       9       E       S       T       `       a       b       l       mL       categories_sizes[$L#L                                                                                                         
              L       default_left[$U#L                                                                                                              L       idiL       left_children[$l#L                      	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c   e   g   i   k   m   o   q   s   u   w   y   {   }����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       Vx�eU��U�8Tٚ�UâU$OT�4CS�;�T�T<��TW�T�fT/ S��UTf8�T�;S*�bTy�dT�lS��S$~�S���T>]^T4S�c�TC�T5tSb�*R͘�T�aJS2c*SxSc�|R��S�YS���R��R���S���S�_HS�S� Q���R�� S<��S���S/�_SѽpSk��SOKT)ÀS�]�Sg�SvZ�S���R�\�R���R�5RS�@S~IPS��ZS��R_��                                                                                                                                                                                                                                                                L       parents[$l#L       ���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <   =   =   >   >L       right_children[$l#L                      
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d   f   h   j   l   n   p   r   t   v   x   z   |   ~����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       B�        BB�RD�` B�  D�  @�ff@��R   A   @�33         D�` D�� D�  D�` B\     B<�H      D�` >���@z�B�     ?�~�   B��Bff   Ap  D�  ?��   A<z�B<�HBa��B4  B�k�   @�j@z�BT��>��j=���A      A�  ?xQ�A0  >49X@���A      B��{@�  ?�/@��B�  Ƥ��D�L����G(qƒf���YZ�1�	F�"GL�DF��G�ݭE��|D��=ƥi�F�4���|L���tJ�ſ�F�j�����&j�(u��B��S�C�ݓ��T2;Ǝ �G�rF	��Ƌ۳En1�G��G{�����uG_aF�wmƃ~�G\��Ž�G"Y'G���H(u�G5��H!F���H
�dGE�c�&�gG�OF�\�G��\�3~�F����/���{���^mG�G5����i9F�9O�?V\��i�F� cL       split_indices[$l#L                                                                                                                                                       
         
                      
                                                                                                                                                                                                                                                                                        L       
split_type[$U#L                                                                                                                      L       sum_hessian[$d#L       F�` FT� E`� E�� F� D�� D�` E� D�� E�( EG  D�� D� D�� DG@ D�� Do� DH@ D�� E_� E� D� D�` C׀ D;� C�  CV  C�  D� C�  C� D�@ C�  D� C�  D@ C<  DH  C�  EM C�  D�� D� D@� D�` D4@ D� CX  CW  C�� C� Cb  B�  B(  C,  C�  B�  C�� B�  B�  C  C{  CL  Ck  DU� B�  CS  C� B�  C�  B�  CY  C�  C5  @�  D+� B�  C�� B  D�  D�  CV  B�  DH� D�@ D  A0  C�  C�  D8� C�  C�  CЀ C�  Ct  C  B�  A`  CI  CF  B�  Cʀ B�  B  CA  B�  @�  B  @�  A`  C  C A�  Bl  AP  C�  A�  BT  B@  @�  B�  C?  B�  CW  B  C!  B,  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       127L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       C�Yp�ݦxG�}���/�i�G�XFH�
ƫ�lF�}��%_Vǚ��G�s�HLn0GV9ƒ�5��$G<׸��
Gn�Ǹ�Y�����=Ǐ�*H+w�G2RHo��G��F���G���߭�~�ƭ#"Ǚd���-mG�h7E�ǁ��F���G�JZ����Ǎ2�+ًF32��.��˧�Ǆ�����*H}lDG�T�G�NY��pH3yGU��G��{Hq]mE�d�H��Hy�ń�JDt�l�W�Ǿg��9���a�1��:Ɨ����*SƆ�CE�W�F�'�ū�Ź�F\|��ٞ�F����HCF6}RG�Ed�����E��M�ǜj�A/#�3�B��ӟGV�Ğ����[�/��Ɣ����HƐ����<m����ҿ�GR�G��F�8�G���G)�dF\2�Fk��m�GL�:G��}��j�F��E�7�G@M7G�uF��F�&�ŧ_^GY);�m��G��G��tG{���˰��NFH��Ʃ�E�n�����F������kƮ�L       
categories[$l#L       [                         	   
                                  	   
                            
                            	   
                     
              
                               	   
                                                     	   
                                      
L       categories_nodes[$l#L                                                  *   ,   -   0   7   ;   >L       categories_segments[$L#L                                           +       ,       /       0       1       3       A       C       D       F       T       U       V       W       X       YL       categories_sizes[$L#L                                                                                                                                                   L       default_left[$U#L                                                                                                               L       idiL       left_children[$l#L                      	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c   e   g   i   k   m   o   q   s   u   w   y   {   }����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       U�`�UU_)nTNp&S�%�U� T7�eT,�@Tf�6ST�XR��@T�y�TKM�S�0S*8�S�լSy�JS�ĳTD:Q��S\ QN!�R�'�S��hT25�S���S�v�Sa��S�R�U�R �Sk�jR#�RV��SSQȫS��?S1n�So�P���QH� SGS�<N� P�A�R�gPP��STx0S��LS�\�R�o�T��R�/�SZ�{R���S(G�R��S�(HS�;Rx��RA4Qρ`QĿD                                                                                                                                                                                                                                                                L       parents[$l#L       ���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <   =   =   >   >L       right_children[$l#L                      
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d   f   h   j   l   n   p   r   t   v   x   z   |   ~����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       B�        D��    B�     B8  A   B  B  @L(�   D�        B   @	��B@  A�     A�R         ?�hB�ffB�  ?�(�   D�@ @b   A�R?A%BP  ?��D@   @&A�  A�  ?xQ�   @���      ?�ff>&�y   @�z�@@  >�VD�` D�@ ?�r�   @IG�@��=ě�   B�(�B�     �a�1��:Ɨ����*SƆ�CE�W�F�'�ū�Ź�F\|��ٞ�F����HCF6}RG�Ed�����E��M�ǜj�A/#�3�B��ӟGV�Ğ����[�/��Ɣ����HƐ����<m����ҿ�GR�G��F�8�G���G)�dF\2�Fk��m�GL�:G��}��j�F��E�7�G@M7G�uF��F�&�ŧ_^GY);�m��G��G��tG{���˰��NFH��Ʃ�E�n�����F������kƮ�L       split_indices[$l#L                                                                  
                                    
                         	                                                                                                                                                                                                                                                                                                                                                L       
split_type[$U#L                                                                                                                  L       sum_hessian[$d#L       F�` F?$ E�8 E�� E�p E"  Ep E� E%� E/` E� D�� Dl� D@ D�@ EiP D� D�� D�  C�� E� C�� E� C�� D�` D.� Cw  D  CЀ D�` C�� EA0 D � CS  C�� Dc� C�� D;@ D#  C  C  EP C�  B�  C^  D�� C�� C  Ck  Dh� C�� D!@ BX  CB  BT  D� B(  C�  B�  Dg� C  B�  C1  EP D7� C�  C�  Bx  C  C�� B8  D� C�  C�  Bd  C  D@ D	@ B�  C  ?�  B�  B,  D�  CT  B,  C�� B�  ?�  A�  CL  D�� C�  CW  B�  B�  B|  C-  Bx  C�� D%@ BX  C�� C`  CҀ AP  B$  C  B�  B   AP  C3  C�� B   @   Cp  Bx  A   B�  DG@ C  C   A�  B�  @�  B�  B�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       127L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       Cm���@��G�ɠF�S���SPH�0G(���&l�GF�#�'�E��2Ha��G���G�@He�!GC�4��G��EF� ��G]�Ɲj����F��H7$H�לG_�KHO�F38G��H���Ǥ#�H.LWF̫Aơ�F~RgG��H1k�D��Gu�m�3��ǔ�Ƹ~G��ǸƷ4�G�m�Ed�H��pG�8�H5�H� �$3G�P�o��H��\Fa|��ų�H�aF� =G�H���G]guȅ�lF�X�G��DC�6LF�����F��FN��G1��F>��Gzl�G��F�[�Ĥ
F�|����XƷr�D�Qƽ��Ɔ��Ŝ:�ƌ);G�,�F� �W�Y��&��ƀ�hG
M�f��F����#Gψ.F�a�F	QG���G���G")����G����5�ǡ��GN(�FL�F��=�ٺG��	G�0�9��Fh������bxG�jG�SEA�MG{�K�	��G�"�GِLƉ�G#{�ƪE�Ƿ�DƵ�GL       
categories[$l#L       7                               	   
                                        	   
                                   	   
                                         	   
            L       categories_nodes[$l#L                   )   -   8   9L       categories_segments[$L#L                                                  (       )L       categories_sizes[$L#L                                          
              L       default_left[$U#L                                                                                                                     L       idiL       left_children[$l#L                      	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c   e   g   i   k   m   o   q   s   u   w   y   {   }����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       U�]�T�F�T�k�TAe�TXZ�T���T��SL��TB�S��SԡS�]@S�$�ToSc�S
 S � S��TSs��S��S��,R��2S�ضT��S��S�S�,hS�S�;�S&hRn�RѬxS(�R��vS �S��fR���RŘS�B�R��`Qc0@S+�fR���Q��R�)�SҎ�So?ES� S�OvR�xSMi@R倍Sw�4R 0S� S�Q��S�2`R�ӎR�ǥS�Q���O�:                                                                                                                                                                                                                                                                 L       parents[$l#L       ���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <   =   =   >   >L       right_children[$l#L                      
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d   f   h   j   l   n   p   r   t   v   x   z   |   ~����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       B�        BM\)D�� @�p�B�  >��@�Q�BW��B,�D�� B�ffD�� @�  D�  D�@ D�@ D��    B�  A�  @��D�� B�  D�  ?a%?�/@��B��C  D�` D�� B�  A33@�R?�#>9XA�@   D�`    =�%>�ȴ>�V   > Ĝ@�  B�  =��=y�#B(  >�n�>��@&>��      B�  >���=�j@�  B�  F�X�G��DC�6LF�����F��FN��G1��F>��Gzl�G��F�[�Ĥ
F�|����XƷr�D�Qƽ��Ɔ��Ŝ:�ƌ);G�,�F� �W�Y��&��ƀ�hG
M�f��F����#Gψ.F�a�F	QG���G���G")����G����5�ǡ��GN(�FL�F��=�ٺG��	G�0�9��Fh������bxG�jG�SEA�MG{�K�	��G�"�GِLƉ�G#{�ƪE�Ƿ�DƵ�GL       split_indices[$l#L                                 
                                                                                       
   
                                                 
                                                                                                                                                                                                                                                                                            L       
split_type[$U#L                                                                                                                               L       sum_hessian[$d#L       F�` Fi� E� E�� F   DR� D�  E(0 D�@ E�  E%� CĀ C�� D�� B�  D  Ep DD@ D�  E�X E=� DQ� D� C�� B�  C�� B�  D{  C�� Bh  A   A�  C�  D�� D  D  C1  DQ  C΀ Em� D;� E7� B�  B�  D3� C�  D�` B�  C  B8  B�  C*  CM  A@  Bx  Do� B8  CF  B�  A`  B0  @�  @@  Ap  A0  C�� C!  DĀ Bl  C�� CI  C,  C�  B�  Bh  BL  DD@ C�  B�  C�  ES  D� C  E C�  A  B�  B�  B  C�  Cb  C�� C  C[  D�  B�  A�  B�  B<  @�  B  @@  B�  C$  @�  B�  B�  @@  A  B  A�  D"  C�  A  B  A�  C2  B�  A@  @�  A   B$  @@  @@  @   @   ?�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       127L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       }CiȐ�{��G�Lőr'���GMUk�D��Di�,67��F��*G*a�H)�F�Bcƞ�#���E�.(�6R4F�|A��n��<�Gw��9�xGyf�F!QH*���vA�G�c�F��d�:`�sJǆ('ƾ�F���7��"fǏ�b��.G�Oƥܜ�j~�@G��Yƫ�H$��F���ǘc�G��Gs�GA�ſ
�H��G�U�G�5��܂H"�5�*��2F�jG6ڇ�Qc#�2ĘF���Ʈ�8���Ѷ+�6m#F��\E�7�Cþ��	Gh���E��G�Ʋt9ƽ�F3mÆ��G�G�����cZ�7!�����3]IƋ��F��G����muRF�?�F�7G���De%G2��O���A�G=F~5�œ�7Fm�gF��GH��DN�bƧ�>Gv@ZF�B�G�s���a��YϹG���G�CF��F�����E�k���{�E0��FY��G b�F���h�EYF��Ƙ��F�q����YL       
categories[$l#L       C                         
                            	   
                                                     	   
                     
                                                          	   
                     L       categories_nodes[$l#L                      	                  !   "   '   )   3   ;   <   =L       categories_segments[$L#L                      
                                                 '       +       ,       -       0       1       2       @       A       BL       categories_sizes[$L#L              
       
                                                                                                                L       default_left[$U#L       }                                                                                                          L       idiL       left_children[$l#L       }               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c   e   g����   i   k   m   o   q   s   u   w   y   {��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       }UF-T)��T�?wS���S��T[��R�AS��wR�@R��S��T�SYhQǔ�R�PR�&pS�/Q�ېR�OR���R�@Ss�bR&ndS��SR�>SahR�zRN��Q�x+R*�rR):�Q�0R�zSY��S3a�Q�PQ��pQ�$�R=ˏRN��RG�`Rz�`Q\F
R0e�R�LhQS�rQ��S� �SNhnS׫S��SM2�    R��<R��Q�8P�v�R �jQr��QG&�R��Q̏ Q��E                                                                                                                                                                                                                                                        L       parents[$l#L       }���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <   =   =   >   >L       right_children[$l#L       }               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d   f   h����   j   l   n   p   r   t   v   x   z   |��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       }Bx           @�ffB�     B�
B�     @E�            A�
=@���A0  ?c�
D�� C
  >Õ�>���   >/�B�  @�  >cS�?�(�=49XB�  Ap  @w
=      =��D�  D�� BQ��   ?�
=   >�-BHD�� A"{?�@��R>	7LD�@ ?�ff   G�U�? A�D�� A   ?&��>�$�A           >�Ʈ�8���Ѷ+�6m#F��\E�7�Cþ��	Gh���E��G�Ʋt9ƽ�F3mÆ��G�G�����cZ�7!�����3]IƋ��F��G����muRF�?�F�7G���De%G2��O���A�G=F~5�œ�7Fm�gF��GH��DN�bƧ�>Gv@ZF�B�G�s���a��YϹG���G�CF��F�����E�k���{�E0��FY��G b�F���h�EYF��Ƙ��F�q����YL       split_indices[$l#L       }                                                                                                                 
                                                                 
                                                                                                                                                                                                                                                                          L       
split_type[$U#L       }                                                                                                           L       sum_hessian[$d#L       }F�` F5� E�X E� Ey@ Ez� D�� EҸ D^� Em CC  Eg@ C�� C�� D�` D]@ E� DV  B  D�� EP B�  B�  E� D�� C�� A�  A�  Cu  DR  C� C�  D� EF` E'� D4� C  A�  A0  D�� Cp  E� AP  B�  BL  A�  B`  D�� D�� C�  Dv� C�� A�  A`  A`  A`  A�  BX  C?  BT  DD� C�  A�  Cz  A�  C�  C�� C�  E(� DҠ Dy� ?�  D4@ ?�  C  A@  A0  @�  @�  C�  D=  C  B�  D�  D�� A@  ?�  BH  A`  A�  A�  A�  @@  A�  B   D� D-  C�� DB@ C�  Bx  DY� B�  C  B�  A  @�  AP  ?�  @�  A   @@  AP  A�  A�  B�  B�  A   B,  D  Cs  Cw  C-  A0  A�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       125L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       }CM���ŦuG2ҡE�#�Ɩ�G��MF����"F�l�EA���ǽ�H��Gy��Fa�G�R�`�mF�]	Ƥ�F��A�MrG�ɢ��QHr��HhjXG�
�H<fKGO�UG�!�Y�G���Z�W���w�VG�E�G�e��t>��r@4G.��F�E����^GS�VH������z�G���G�&H���B<��	�qH�jHk�r�g%��:cOG���HE�zF��_Ƶu�G��G�f�H�|�ǽYUG�;����]���?C�SL�F?�x�DP�G0?�$�E�%*�����SJ����GD	FAoE�(��d�lEn�,����G��GS��R�GsGřE����
�&�l>NEF���E>�jutG.�(�&�dG�1vFg��"�����G#���jSGU�$G����7�G,���E��E���#�`Fŕ��7��F^G�͸Fp��7���c���ҤGk��D3�G	�����Hg��>��7���jǮG#���.�L       
categories[$l#L       ?                                       	   
                                          	   
                                  
                                
                           	   
               L       categories_nodes[$l#L                               "   #   '   +   ,   9   =L       categories_segments[$L#L                                                                       )       *       +       0       ;       =L       categories_sizes[$L#L                                                               
                                          L       default_left[$U#L       }                                                                                                               L       idiL       left_children[$l#L       }               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [����   ]   _   a   c   e   g   i   k   m   o   q   s   u   w   y   {��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       }T���T)�S���S�p�Sw
hS��4S=OR�.5S�T3Sq��SRJ<S+h�Sna�S)��SxR�R�R��XR8|S|ȬR���S6b{R߅�R�xS6�S:,S%��Sz��SɭS
P�SLМR�Q��R�	lQ�iRmh,Qʹ�QZE S7R�:R��R��Rx֨Rl� Ra�@R�Y�PÑd    SXHQ��gR��/R�jpSPՄRi�^S�(Sm�HR��rS �R�s�R޶�R�Z�R�~�Q�:�Qs2/                                                                                                                                                                                                                                                        L       parents[$l#L       }���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <   =   =   >   >L       right_children[$l#L       }               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X   Z   \����   ^   `   b   d   f   h   j   l   n   p   r   t   v   x   z   |��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       }B�33      B@        B�  B4     B�  A�  >ؓuD�@    >D�� B#
=>���>{�m@0A�Bh  @@  ?�>>���   D�� <�`B@�
=>ٙ�AAD��D�  D��       @��D� ?��   ?�9X?���B�        B\)G�&=��B�(�>���>���@�  =t�>���?�9XB��B     >��@�\)C     @@  ���]���?C�SL�F?�x�DP�G0?�$�E�%*�����SJ����GD	FAoE�(��d�lEn�,����G��GS��R�GsGřE����
�&�l>NEF���E>�jutG.�(�&�dG�1vFg��"�����G#���jSGU�$G����7�G,���E��E���#�`Fŕ��7��F^G�͸Fp��7���c���ҤGk��D3�G	�����Hg��>��7���jǮG#���.�L       split_indices[$l#L       }                                     
                                                                              
                                                      	                	                                                                                                                                                                                                                                                                     L       
split_type[$U#L       }                                                                                                               L       sum_hessian[$d#L       }F�` Fk E� E�P E�� De@ D�� EN  E�@ DΠ E�0 C+  D:� D�@ C4  E;@ C�  D/� EZ� D�  B�  E�� A0  B�  B�  B`  D,� C�  D� C  A�  D�� DϠ CO  B�  D� B�  D�� Dɀ D�� C�  BH  A�  EK` E$P @�  @�  Bh  A   A�  B�  B<  A  B�  D� A�  Cـ D
� B@  C  A   A�  @�  D�� A�  D�` C2  B�  C
  B�  A�  B�  D  Bp  A�  BH  D� D�  C  D�  C]  C�  A   A�  A�  A�  @@  E  D5  C�  E� ?�  @�  @�  BT  @�  @�  A�  A   A  B�  B  A  @@  @�  BT  B  D� B�  A   AP  C�  B�  C�  B�  A�  A�  B�  B  @�  @   Ap  @�  @�  @@  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       125L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       C;F����]�E>rG&� ƖnA�?�G�8�F��G�R�E�
��$'������QG�Y0Fo�+G��F��7Ɵ0�Gv��H-�NF�ZC�d�U-��j�ƭoſ��F�+���g&F��iH
��G�J+E��G�R��́�G1��� [ư�Gt�MH��HGeC�G�#HT��ƍ�|G7��}0�H�=Ǜ��/YR�DN���~E�I�ȸ�ƚP|E��F��NHn��P	G"�G�+�Ǫ_4HeW���Gw1EyM�G��D�qHF��vGp*����F�%łq�F��$F��6�U��ůKP��� � �KG;��Fp�bH�HF��TFTG]���H��G<� G��3�ݤ-GE �FB�Gw>e�졑�y�D� G��_FQh���C#�cD�E�%�ŋ[0Ǝ,Eż���A���Ž�F9�XF��v��u��T�EhE��8ŗ��ExU^F�{wG�oŤ1��~eYE��zG	�e�c��G�eF�[F�����}GUT'��U��WVM�f��L       
categories[$l#L       "                            	   
                                           
                   
               L       categories_nodes[$l#L       	                .   2   6   8   >L       categories_segments[$L#L       	                                                                 !L       categories_sizes[$L#L       	                                                 	              L       default_left[$U#L                                                                                                                     L       idi	L       left_children[$l#L                      	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c   e   g   i   k   m   o   q   s   u   w   y   {   }����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       T ��T	;�Sg�>S�;"T-^�R�((SO�KS�˧S$��S���Sy�Q(S�R���S�	R���R��(SE3�R�SER���S�؎SPp�Sa��R��LQ#P� Rq�RyShR��|R��zS/OR��tR��RQ��S#b�S�hR�5RFYS'��R�=�R�N�S8�R��SR8R���R�#$RQ��Q��LQ��P���Q� P�ېQ��TRژQ>UpRuj�Rn�Q�nR�XES�9�S�
RC!LR~>�N�                                                                                                                                                                                                                                                                 L       parents[$l#L       ���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <   =   =   >   >L       right_children[$l#L                      
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d   f   h   j   l   n   p   r   t   v   x   z   |   ~����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L          D�� BNG�D�  @�
=B   B�  B�\@/\)B��=D�� A�=q@�     ?��D�� @�     B�ff=���>^5?@�  @�  @�  >,1   D�� A@  @�ff>���>��/>p��?��B�  >cS�>Y�=oB��>y�#>�J@�  =��`@�  A�  B�  @�     D�` ?!G�D��    A�  <D��A�     D��    ?�@E�B�  Bn  =�j   Gw1EyM�G��D�qHF��vGp*����F�%łq�F��$F��6�U��ůKP��� � �KG;��Fp�bH�HF��TFTG]���H��G<� G��3�ݤ-GE �FB�Gw>e�졑�y�D� G��_FQh���C#�cD�E�%�ŋ[0Ǝ,Eż���A���Ž�F9�XF��v��u��T�EhE��8ŗ��ExU^F�{wG�oŤ1��~eYE��zG	�e�c��G�eF�[F�����}GUT'��U��WVM�f��L       split_indices[$l#L                                                                       
                                          	                     
                     	                                                                                                                                                                                                                                                                                                             L       
split_type[$U#L                                                                                                                             L       sum_hessian[$d#L       F�` E�  F+@ Exp E� E�� E�� D�@ E/� D�` D�� D  E�X E� C  DL  C�  D@ E� Dj� C   Dp� CK  CD  C�  E:� DӠ DT  E�� B�  B�  B�  D2� C�  B�  Cz  C�� E
� Bd  A@  Dg� B  B�  C�� D� CH  @@  BT  C  B�  C�  C�  E#@ DB� Dd� DR� @�  E�� C�  BH  A�  B|  @@  B<  BX  A�  D.@ CJ  B�  A�  B,  B�  C#  A�  C�� E  B�  A�  A�  @@  A  C�  D� A@  A�  B�  B  C�� A   D@ A�  B�  B�  ?�  @   @   BL  C  A   A�  B�  C  C   C�� B|  A�  E" C�  C�� D� C�� D(� C'  @�  ?�  En� D� C  B�  A0  B  @�  A�  B`  @�  @   ?�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       127L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       yC7�Ez K�������F�M�ƿ�0�QuD��VƠ�cG:�E�3aƍQ��eR����R�F&�.��`m�*���+�G���F�BF��k�_ە�3����u-�	��F�U�H <��0\SGL����vFk�d���O�-7E����]3tGD)�`an�зX�0�{G��G
$]Ǹ��E�d$G�E ;��.cBž8��oy��w�΢�� ��ǲ��ƭ?<G�EFG�L�ŔJU�X�(G-��F�^@�<�gG� ��hD�3,FE:��M}F֋����/�jFY��`���y��2	.G+DEQ�9�����E�\�J=eF��Wǒt(G�u� ��GX��FƍGeN��9H�D��"G��\G:�{E:8E��$�7���x9�F������2�S�ͻ�ƒ����}ƀG#��1E!�4�ge������:��h�E������E)�qGBmtF=��^nzŽ��ƿ��G\��F�Tþ�g�-bJ�<�L       
categories[$l#L       R                                	   
                                   	   
                         
                	   
         
                               	   
                             	   
                               	   
                        
      L       categories_nodes[$l#L                                      "   ,   /   8L       categories_segments[$L#L                                                         %       (       5       6       @       L       QL       categories_sizes[$L#L                                                                             
                     L       default_left[$U#L       y                                                                                                      L       idi
L       left_children[$l#L       y               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c   e   g   i   k   m����   o   q   s��������   u   w����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       yS׫ZS�\R*-(S:��S�նQ�	pRO;8S6S�R��rS�l�R�RQ�j�Q��Rk�4Q�� SJ��Rt`rR�
$Q���SMv�S��SMբR���Q�
�Q1�Q���Qˉ�Q��(R-+|PPH(Q��hS{UCS)E�R9�R���RS��R���R �`R3�S�k�S_pS~��S;�*R�`�S��RXcR���Q�ϊQ�4Q)D�P��Q��XP��Q���QUJB    O�*nR�RI�        O��P�1�                                                                                                                                                                                                                                        L       parents[$l#L       y���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   8   8   9   9   :   :   =   =   >   >L       right_children[$l#L       y               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d   f   h   j   l   n����   p   r   t��������   v   x����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       y   B�ffB�\?��      @���      @L(�>��F@�  B�  @   >1'?�V>�7L@kC�?�9X=��B0  >�"�   @�  B�     >?|�   C     =]/D�� ?��B�   @�Q�@o�w?DZ?��D�� CW
D� =��A�     ?��A@     Bg��B���D�  >.{>&�y=�oB0  G�L�   =ě�?У�F�^@�<�gB��@�  D�3,FE:��M}F֋����/�jFY��`���y��2	.G+DEQ�9�����E�\�J=eF��Wǒt(G�u� ��GX��FƍGeN��9H�D��"G��\G:�{E:8E��$�7���x9�F������2�S�ͻ�ƒ����}ƀG#��1E!�4�ge������:��h�E������E)�qGBmtF=��^nzŽ��ƿ��G\��F�Tþ�g�-bJ�<�L       split_indices[$l#L       y                                                   
      
                                                	             
                  	                             	                                                                                                                                                                                                                                                                             L       
split_type[$U#L       y                                                                                                            L       sum_hessian[$d#L       yF�` Fl� E   F6� EWP D� Cu  F� D�� D�� D�� D�` D@� CI  B0  E�@ E�� D�� D� C�  D�� D�  D)� D @ C�  D9  A�  @�  CD  @@  B$  E�  C�  Es� D�` D�� B�  C�  C~  B$  CĀ D�� B$  D�  B�  C�  Cr  C�  C  C�� @�  D2@ A�  A�  A  @@  @   C0  A�  @   ?�  @   B  EG0 D�� C΀ B,  DJ  EAp Cڀ D� D�� C�� A�  BD  CN  B�  B�  C;  A�  A�  C�� A@  B8  D�� @�  B  D~� @�  B�  BD  C�� B�  Cf  A@  C�� Bl  B�  B   C�  BL  @�  ?�  C`  C� @�  A�  A`  @�  @�  @�  ?�  ?�  B�  B�  A`  @�  ?�  ?�  B  @�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       121L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       }C^mF�!�?|sG$�HFŏ��G.�G��F�CF�2�� ��E�[���\F���G��)FAגG�����QGQJG���%��Q�G�eF�g>��@��Y�%�xFڢ�ǋ�<H>�É�E.�FG~w�H�g�G�}�Ge1�Ư�G��H��o��GP��E�@[�!�L�^�DQ�H"߽E�wUE螬Ga��F�zH�'d�4]4E�J\�c�DǍ�Fk,TGݬ<ƕ�ǝ8NGӭ�Hɸ��Q�>F����*BWF��uƦKF�1�F�FH�G`�F�dF˴���EG2�ƕ��B+3 F�MIG��"F&��G���+n�F�ezE��É�FF�Ǖ����/��@cƮ����R�E�ZFp��G���E�4š�F	�G���E�7�Gf.F�a�Əs^��Io�����}���F��D�eRF�Ə>Zƃ���hBFH�gG�GVl9���F"C���)G���F�BH_YF�E�ǭd�Ɛ�@����F�BL       
categories[$l#L       F                                	   
                                  
                               	   
                                              
                                  	   
                              L       categories_nodes[$l#L                 	            +   .   3   4   5   8L       categories_segments[$L#L                                           $       &       )       *       +       2       @       EL       categories_sizes[$L#L                                                                                           L       default_left[$U#L       }                                                                                                        L       idiL       left_children[$l#L       }               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c   e   g   i   k   m   o   q   s����   u   w   y   {��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       }S|�S�S?͓R�J�R<�dS� S+ES=R���R�s�Q�mxS'%fRÞNR���S�Q�+0R���R���Rd�*R�� Q���Q��}Q�ZS^�R;�HR���R��<R�>�R���S4�ZR~t�Q�MQ�kLR�^@R��QةRv�nR��RR�RP�~R���P�i%R	v�Q<�Q�_P� �N��S;XS��OR��eR�R� �R��R���Q��`R�R���RBo    S'5R<n�Q#��R�L                                                                                                                                                                                                                                                        L       parents[$l#L       }���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   ;   ;   <   <   =   =   >   >L       right_children[$l#L       }               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d   f   h   j   l   n   p   r   t����   v   x   z   |��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       }      B�  @��H?;d>hsD�` BA��?�   AP     D�  @0A�>���>�b@@  >)��B�  =�`B   @   >�S�>���>�ffD�  @-?�/   ?*~�>��A  B��>���=m�h@?��D>��R>߾w=C�@J=qD�� @@     D�` B=�H   >��wB|ff>��HAp           @�  D��    @Ϯǝ8NB�  ?��FD�� ?ȴ�*BWF��uƦKF�1�F�FH�G`�F�dF˴���EG2�ƕ��B+3 F�MIG��"F&��G���+n�F�ezE��É�FF�Ǖ����/��@cƮ����R�E�ZFp��G���E�4š�F	�G���E�7�Gf.F�a�Əs^��Io�����}���F��D�eRF�Ə>Zƃ���hBFH�gG�GVl9���F"C���)G���F�BH_YF�E�ǭd�Ɛ�@����F�BL       split_indices[$l#L       }                
            	                                                            	       	                     
                                   
                                                 
                                                                                                                                                                                                                                                        L       
split_type[$U#L       }                                                                                                                 L       sum_hessian[$d#L       }F�` E  Fg@ DH@ D�� F]� D  C�  CÀ D!� Dn  E� Fh C�� B�  C(  Cr  C~  C	  C�  C�� Dl� @�  E� EP F� C�  C�  B<  B�  B4  C  A�  A`  Cd  Bx  C@  B�  A�  B�  C�� Ch  B  B\  D^� @�  @   D�  C� B�  D�� E�� D�� C?  C/  C�  B`  B  A  Bt  A  @�  B$  B�  A�  @�  A�  A   @�  A�  CJ  B,  A�  B�  B�  B|  BT  A0  A   A  B�  CM  B�  CE  B  @   B  B  A�  D%� Cd  @   @   ?�  ?�  D>� D�� C�� C  B�  A�  D�� C�� E�P D΀ B�  DԠ B�  B�  C  B(  C�  B�  B  A�  A�  Ap  A   BT  @�  @   @   @   @�  B  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       125L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       qB����.E���7���u�E�Yƌ���	BiGp�5�	~�GV0F��D�H��Uj��۝�	)�u��F���E�g�����RYFX�G�ܜG&�2E�h��O��G\�B�;b��]w�D��~�Qm��;��瀌Fy��q�����G��N�5�sG��nŏ]G��HGolH&�6G��gG� Eo"H$m����JF �H>{�G!B��C#�G� Eޮ&ǹ�Ƨ$uG1g���ӃǏ�����ѻ�h����Ā��F��I��d�ƲfĊ�<�n��Œ{F��D��ƜOF���g4E�q��!��G����omE���Gz|�G^W�FJ�aD��G'!]�ܟ�F��E<��.�GS&�Ɔ��7�=F-	��G�Fcp���5G�� E�}G1ŕ(�E�,*F�;4Ţ:6�.R}Ɩ��D���Ʋ@�F��|�GӇƒdFa�)������L       
categories[$l#L       1                                   	   
                        
                                   	   
                                                      L       categories_nodes[$l#L                            "   #   *   6   7   :L       categories_segments[$L#L                                                  $       +       ,       -       .       /       0L       categories_sizes[$L#L                                                                                           L       default_left[$U#L       q                                                                                             L       idiL       left_children[$l#L       q               	                                    !��������   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c����   e   g   i   k   m   o������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       qS2ؿR�n~S=��Q(I(RQ�|SE�:Q�)�P߀�Oe0RY�RRmSw��S
Q��bRy�P�� P�2F        Q�PR8R��Q�8SphS�R�>XR�E�R�4Q���Q��R,�vP�P�Q�(P��HN�� Q�|P��DR׺Pp8�Q�)"Q���Qz(�P�mPS6�S�8R���Q��HR���S
	�R��R�p�Q��@    P��QKTQw�Q���R{R�D                                                                                                                                                                                                                        L       parents[$l#L       q���                                                           	   	   
   
                                                                                                                             !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   5   5   6   6   7   7   8   8   9   9   :   :L       right_children[$l#L       q               
                                     "��������   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d����   f   h   j   l   n   p������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       qB5\)A�
=   ?��FB�     B�\A  @@  A"{>�ƨ@�z�A@  A     >(��   F���E�gA�  ?���=��D�� D� ?�9XD��    A?�M�@,(�>�`B   @�  A�        A�  ?�M�@�  =m�hB-��B0�\   >�bD�� A,��?�p�Bp  ?   @   ?�oD�@ G� @@        @6��B��   ����ѻ�h����Ā��F��I��d�ƲfĊ�<�n��Œ{F��D��ƜOF���g4E�q��!��G����omE���Gz|�G^W�FJ�aD��G'!]�ܟ�F��E<��.�GS&�Ɔ��7�=F-	��G�Fcp���5G�� E�}G1ŕ(�E�,*F�;4Ţ:6�.R}Ɩ��D���Ʋ@�F��|�GӇƒdFa�)������L       split_indices[$l#L       q                                  	                                                                                                                 	            
                                                                                                                                                                                                                                                  L       
split_type[$U#L       q                                                                                                     L       sum_hessian[$d#L       qF�` E�� F9| C؀ E�  F#� D�� Cր @�  E� B�  EO� E�H D�  Cu  C�  A�  @   @   E�  C"  B�  A�  D�  D�  Eؘ CV  D�� B(  B�  C1  C&  Cj  A�  @�  E�� AP  C  A@  B�  Ap  A�  A@  C)  D�� D�  A�  Etp E<� A�  CB  D�� ?�  A�  A�  B4  A�  B@  C  B  C  B�  C%  A�  @�  @   @@  Ep E
� @   A0  B,  B�  A0  ?�  B,  B  A`  ?�  A�  ?�  A   @   BH  B�  D� D"@ D�@ Cw  A�  ?�  EdP C�  D�@ Dt� @@  A�  C   B  Dw� B�  @�  A@  A   A�  A�  A`  A�  @�  A�  A�  B<  B�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       113L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       wB���D�|��ϙ�:�F�sƤ:1�WV1ƌ��Ğ��E<�F�����j���@�.��ǎƠ&|�C8jDN.�fV<÷��G�F 1%GR
/Ƽ���ru-�Lq�=��D��G�@ǚ��G{�ƥU�G'��GW��t`F-�\��pCƁ��F�+\F�#Ŏ:PF���H���F�c���/G:�XH9��G����.�`I4E'�ƫjnG���t|Ƿ��E�k�ǘ9�G/r�Fd�bǅ���mk�ƌ
mGC$���š�E*HFֻBF�h\Ƌϳ��C4�E�wÃ���6
'F�\�Y���\EK��F�׆E���G5��@�,F� 6ĮpE�EG���G�|E����
w�#�F�&QE_�9H}F�:F���T�tF.N�,��E�5�ƣ���T6E�C elƃO�H��F	A��Qd�E���	�o�mfż�DFz��߸�� �F����p�ݒ�L       
categories[$l#L       $         
                  
                          
                          	   
                              L       categories_nodes[$l#L                         #   ;L       categories_segments[$L#L                             
                            L       categories_sizes[$L#L                                                        L       default_left[$U#L       w                                                                                                       L       idiL       left_children[$l#L       w               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c   e   g   i   k   m   o   q����   s   u��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       wS US �QؠXR�JS-��Q���Q��HQTpRz��R�%(S�Q
Q���Q�uRQe��Q/xQRT�R]�iQ���R���R�uR�/NR�XQGȲP�kdR# �Q��8P��Q"	�Q�	\Q<�<Q6�PiW~QlDP�RG�'R��Qm8(Qx�R���R�;JR��`QG`@R�R/Q�=�R���S��P�5xP�+�PP��QީR�Y�Q�U0Q�PO��P    P&� Q�.�                                                                                                                                                                                                                                            L       parents[$l#L       w���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   :   :   ;   ;L       right_children[$l#L       w               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d   f   h   j   l   n   p   r����   t   v��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       w?�ffBo33D�� Bff?"J   B4z�B,     Bp  D�  ?�@bN@c�FB�  ?�G�B8  @	��A@     >�$�   B�     D�` B�  B�\?��@��B�(�?wK�>��@�B z�=H�9   ?�9X>��!BNG�A�  =��->]/B�=q=#�
?��?ȴ9B�ff@��>O�=�l�?��H@@  ?�Brff@c�FB�
A�G/r�@kC�   �mk�ƌ
mGC$���š�E*HFֻBF�h\Ƌϳ��C4�E�wÃ���6
'F�\�Y���\EK��F�׆E���G5��@�,F� 6ĮpE�EG���G�|E����
w�#�F�&QE_�9H}F�:F���T�tF.N�,��E�5�ƣ���T6E�C elƃO�H��F	A��Qd�E���	�o�mfż�DFz��߸�� �F����p�ݒ�L       split_indices[$l#L       w                                                                                                	                                  	      	   	   
      
   	                               
                                                                                                                                                                                                                                                L       
split_type[$U#L       w                                                                                                                L       sum_hessian[$d#L       wF�` F�� D9  F&  E�` D@ B�  D�  F  E�0 D�� C�� C�  B  B�  Di� C  F � D�` E�  C�  D3� D� B�  C7  C&  C,  A�  Ap  B�  @�  Dg@ A  A`  C  D�  E�� D�` B`  D� EX� C�  @�  D� B�  D� A�  A0  B�  A   C/  C  A0  C  B   @�  AP  @   AP  B�  @�  @   @   C�  D#� @�  @@  A0  @@  B   B�  Dn� DI� E�P BL  DO� Cƀ B,  AP  D� Ap  C�  EB  Co  C1  ?�  @�  @   D@ B�  A   C�  CG  @�  A�  @�  @�  @�  B�  ?�  @�  B�  B�  B�  Bt  ?�  A   B�  A�  A�  Ap  @�  @@  A  @�  A   @@  B   B,  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       119L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       [B��Ei��%�(D�:UG*��)��G�\E��@�
�F��2H�^����Ԕ8ık�F3�&���HƦ�F���Ǵ^SGL�Hr��ģV*�O��F[ƟB5ē���Q�nFa���u��.ŋ������_5�F˚dG�[_�]	Ƹ�|D��G\��FʤH�xGB�c�>�V�5���y4 �1DCF���Ƅ��th�Ei���I������[WE�H�D�����aƧ�|�ɽX�^(v�ر.�����ƛ�B�6V���FK��/�Jąw�ǚ�F��d�`���InF��F�> �i��F��TG��\G���D֩r�e�{ī�����ƌ}�c�F���G0 E�h��K�EW���p�FE�eL       
categories[$l#L       2               
                    	                               	   
                  	      
                                               	   
            L       categories_nodes[$l#L             
                  #   )   +   .L       categories_segments[$L#L                                                                       !       "       $L       categories_sizes[$L#L                                                                                    L       default_left[$U#L       [                                                                              L       idiL       left_children[$l#L       [               	   ����                                 !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A����   C   E   G����   I   K   M   O   Q����   S   U   W   Y������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       [R�E�R�c�Rn[�R��_S��Rkj�    R�IQ�z�R��R��R�I�R��%R�̱S>Q��Q��R���R/,R>UPRP�QΉ�R���Rb�@R2��R��R�"R�8�R��~Q5p0Q�?�Q��QP/yR���    QP�`RB�R��    P�^[P���Rz�Q*�lQ��    R
�SR�c�R1$Rx\                                                                                                                                                                        L       parents[$l#L       [���                                                     	   	   
   
                                                                                                                                         !   !   #   #   $   $   %   %   '   '   (   (   )   )   *   *   +   +   -   -   .   .   /   /   0   0L       right_children[$l#L       [               
   ����                                  "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B����   D   F   H����   J   L   N   P   R����   T   V   X   Z������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       [@.v�B�ffA�     >�33@���G�\D�  D�� ?�r�      @�\)@�  @
=D�� ?J~�?���>���A   >z�>D��B�  @�   @@  >D��      B-��   D�  @E�?��`G�[_   @�  B�  G\��@   ='�   D��    �y4 B�     ?��D?q&�Ei���I������[WE�H�D�����aƧ�|�ɽX�^(v�ر.�����ƛ�B�6V���FK��/�Jąw�ǚ�F��d�`���InF��F�> �i��F��TG��\G���D֩r�e�{ī�����ƌ}�c�F���G0 E�h��K�EW���p�FE�eL       split_indices[$l#L       [                	                                
      
                                                       
                                                	                                                                                                                                                                           L       
split_type[$U#L       [                                                                                L       sum_hessian[$d#L       [F�` F^\ E9� FY� C�  E9� ?�  F-4 E2� Ci  BL  C� E� EĀ E�� E� D � CU  A�  A�  A�  CE  C�  D�� D�` E�P @�  E�X C�  C  E
� CQ  C�  CQ  @�  @�  A`  A�  @�  @�  A�  B  C#  C�  A   D?� C�� D�  B�  E E�H @@  @@  E� E� C  B�  B   B�  D�� C�� C5  A�  C�  A�  CI  A   ?�  @�  A   @�  @�  A`  @   @   ?�  A�  @�  A�  A�  C  B�  C'  D:� A�  BX  C�� D� Cj  B�  A�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       91L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       B���Eo��Ť�7�	�FI�2F<���� ��P6��**�FSFGy��ҘgF�K��u��>�eE&�y�Z�	ǥt6ơ�>FX���O=/G�#�Fת�+8�G�.GT�����G���Ƃ��E���:i}E��M�*�ƅ�G~r�GoV0ǲ����F�U{F�0DD����Î9�X�9FB3>Hal�U��G��H�!��ǁ�-G3�H	2F\��GĢpE�a�π	H%���
*Pƿ���˰�E���HsU��O�Y�D�p<G-@���(C��ť�>G���G�uGu89Fͅ��#�Ƭ.��"������+�F�:.��}-E��F���E83)��C�$z�F3���rZ����GJŠzQF�yG����=�����,Gp&�F��BF���H�5���F;<�FGv�ę�F��qG\uā��FL�G�s�jj#�*gFL��NN�E2^G�ۭE�<PE8v��/ş���Q=}D��+ũ�6D��Ƙ��F=
G�o�SF7[jƚ�SG^��L       
categories[$l#L       9                     
                             	   
                              	   
                   	                                      	   
                        
         L       categories_nodes[$l#L                    	            #   (   *   1   7   8   :L       categories_segments[$L#L                                                                              "       #       $       1       2L       categories_sizes[$L#L                                                 
                                                        L       default_left[$U#L                                                                                                                 L       idiL       left_children[$l#L                      	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c   e   g   i   k   m   o   q   s   u   w   y   {   }����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       R��ZS �R��mR�.�S8�R�ýRZ��RV��Rr�R�?�R�RRY�R��1Rw
|RqE�R��cR_�wQ�D�Q��0R�h�R ��R��R�#�R;�rQ� R�QS�RO�R0lR�#�R*/R�>RM�(R5p�S��PAN�Q��xQ���Q��BR�^R��QR�R�TQ��RhHpQ���Q�"�R;��R��`N���P���Q�� RY?Q/�"Q �,Q�DQ�1R<�(R�R`�#Q'p0R�8Rf�j                                                                                                                                                                                                                                                                L       parents[$l#L       ���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <   =   =   >   >L       right_children[$l#L                      
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d   f   h   j   l   n   p   r   t   v   x   z   |   ~����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L          A�     A"{A��>���?)��   ?�$�   A�HA�     <o   @�A33   ?DZ@Z=qB�ff?)��A�  B��=A�  BW��?��>��B   C  D�� @�  ?ߝ�A�  D��    B�  B�  ?�ffB�\   @�   =� �>���Btp�=�1D�  B�     A�  A0  ?��
B��3?xQ�      Bg��   A<z�B{D�� B�  D�p<G-@���(C��ť�>G���G�uGu89Fͅ��#�Ƭ.��"������+�F�:.��}-E��F���E83)��C�$z�F3���rZ����GJŠzQF�yG����=�����,Gp&�F��BF���H�5���F;<�FGv�ę�F��qG\uā��FL�G�s�jj#�*gFL��NN�E2^G�ۭE�<PE8v��/ş���Q=}D��+ũ�6D��Ƙ��F=
G�o�SF7[jƚ�SG^��L       split_indices[$l#L                                   
                                                                                                             	         	                                                                                                                                                                                                                                                                                                                    L       
split_type[$U#L                                                                                                                        L       sum_hessian[$d#L       F�` F� E�  E�� E{� Dq� E�� E� C�� El� Cp  C�  D� E� Ej  E�� Dz  B�  C3  EH D� B�  C  C�  A`  C�  Cp  A�  EP D�` Dڠ Ea  D�` Dq  B  @�  B�  C  B,  D�� D�� C�� B�  A�  B�  B0  B�  C�  B`  @�  A  C  C  C-  B�  AP  A   D�@ D�` D�� @�  D�` B�  E_� A�  D� D#@ Dp� ?�  A�  Ap  @@  ?�  B�  A�  B�  A  A�  A�  D�� C�  D�  C�� C� A�  B  B@  @�  A�  B�  A`  A�  A�  @�  B�  B$  C�� B  A�  @�  ?�  @@  @�  B�  B\  B�  A  C  A�  B4  A�  A  @�  @�  @   Du@ C�� C�� D  D�� B@  ?�  @@  D�` B`  B�  @@  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       127L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       kB�fD5?�ƥC��zчE��^F+��P�ţG=F�;ŜsZE���UՇG1f$�&7��%:�7��Ɲ۟Gʶ�EJ��U���C�F7�&ŦO�~CǸ�QH(?�E�{��6��FE����^G�.-E9�4����D"u�{rIDH�UH�}G�k]��O^FI�Y��5ǉ�.GR�G0�E�.uD�)	�Ղ��k�Ƿ���Ud�Hy��G$2�x
l�����T�y�˴��Q߸EcE����2����6��DiXǁ��_���C�F?�FW@CGxߣFB
G���L��GA�>�}�?F@���:K��ł���	�5G�<�WDE�iG	�]E�T�(�E3ţ�fF���O �D�#:��,�+�őgD�	Z�l�G�j�G6;F��G�K�/����ƃS�ǅ������F�}���s%���ZL       
categories[$l#L       ,             
                         	   
                                             	   
                                 	                L       categories_nodes[$l#L                                  1   6   7L       categories_segments[$L#L                                                                 #       )       *       +L       categories_sizes[$L#L                                                                                    L       default_left[$U#L       k                                                                                              L       idiL       left_children[$l#L       k               	                                    !   #   %   '   )   +   -   /����   1   3   5����   7����   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c����   e   g   i��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       kRZ��R�U�RLJR:7�R�%�R�1�R���RakHR��{R��R�n'RG�R��/Qt?�R���Rl/4R��R��R@�oR*�R%s�S6O R�d�Q�3�    R���R3�ZP��0    R0d    Q��IQ���Q�w�R��LQ�S�R_�TR�5REM<R>w&RJ�R'O(R� SO<`R~�&R	iR*�O��bP�_�Qb��Q��PQ+~�P�x    O�a�R<�R 8                                                                                                                                                                                                        L       parents[$l#L       k���                                                           	   	   
   
                                                                                                                       !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   6   6   7   7   8   8L       right_children[$l#L       k               
                                     "   $   &   (   *   ,   .   0����   2   4   6����   8����   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d����   f   h   j��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       kD�     @�  D�  D�  >���>�+      @�  ?܋DB�  > Ĝ   Ap  @�  B�=q   =�9X=�1C        ?�dZǸ�Q=�\)   BH  FE��?��G�.-D�@ B���A�  >J>�x�@@  B���@�  BrffB�  D�� >~��@��AR{@�  D�� B�  ?�$�   ?hs@:�\B"  ����      BZ  EcE����2����6��DiXǁ��_���C�F?�FW@CGxߣFB
G���L��GA�>�}�?F@���:K��ł���	�5G�<�WDE�iG	�]E�T�(�E3ţ�fF���O �D�#:��,�+�őgD�	Z�l�G�j�G6;F��G�K�/����ƃS�ǅ������F�}���s%���ZL       split_indices[$l#L       k                     
              
                                                                                                      	                  
          
                                                                                                                                                                                                                        L       
split_type[$U#L       k                                                                                                L       sum_hessian[$d#L       kF�` F�p C�  E�p F( C  C�� E�P C�  E@ E�0 BL  B�  Ap  C�  E� Di� Bl  C�� E@ B�  E�x D�� BD  @   A�  B�  A`  ?�  C�� ?�  EO� E0P DG� C	  A�  B  B  C�� D� D�� B�  AP  D@ E�0 D�� C�  B   A�  @�  A�  BL  A�  @�  A   C)  C*  D�@ E@ E  D	@ C�  C�  A@  B�  @�  Ap  A`  A�  B  @�  C�� @�  C�  C,  D�` A0  A�  B  A   @@  C�  C  E�� A0  Dv� C�� A   C~  A�  A  AP  @�  @�  ?�  @�  A  B8  @�  A   A�  ?�  A  C  B  B�  B�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       107L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       }BdT�E������F_��ŚW�E�ŏF��ŵ#�Fb����ń}ǀ�9F7���0[F-�4Gf�'īG��Š݄G$��Ƅ�BEɄ��EL�&���']ǹ��Fd�b���FXM��7��Gp�F �yG�E�����K��j7oHl9��l�sE����@�Ƥ�+G��c�8���M�7G��]�	`.ő6F�x��9/�G���Ǜ���e�F��U���EL�F�r�Ʋ����~BG�D�E���Fs��ƌ��G��ÿ��Ef}ţ+�G?}FP�iF��*ƀ�nE^���ƫ�]G?��G-��G�b7F
�QƯ3G��DK�|��}�A��ňV�	��F�VD5�$C}��ݦ�ŀo3��¼�"FG$եƵ9qD{UX�{������D?�5F�@��@a)�B�GG�)�/�������ǘ%ƅY�f�Ƹ$��=�CȰoF��F�quE�� �	�wF�&*Ʀد�Tp�G0O���pD=qF�19ř��F���Ųj�F�hL       
categories[$l#L       :                          	   
                           
                                    	   
                              
                   	                                        L       categories_nodes[$l#L                                "   #   &   *   +   ,   /   8   ;L       categories_segments[$L#L                                                         !       "       #       '       (       /       4       7       8       9L       categories_sizes[$L#L                                                                                                                       L       default_left[$U#L       }                                                                                                         L       idiL       left_children[$l#L       }               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c   e   g   i����   k   m   o   q   s   u   w   y   {��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       }RC8�R���R� |R��+RA�'R�%�R�"�S�Rm1�R�q�R�R�ԐQ�-R���Q���R��R��R���SP]R�SR�R�%R��sRԟbR�&P�RPQ��R�B4Q�M~R#^�R% ,R\8TQ� �R��(Q��JR,;-R��R.LQ�/Q�N�RY�Ql�R���Q���RV��R~`�R#�9Rd�GS�|R#�QCjdP�Z�P�\    QTg�R0gR�FlQ���P��HQʦQiR��!QͦZ                                                                                                                                                                                                                                                        L       parents[$l#L       }���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <   =   =   >   >L       right_children[$l#L       }               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d   f   h   j����   l   n   p   r   t   v   x   z   |��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       }>� �   ?"J?���>z�?S��?)x�B�B�?�? �@P  A�D�� @�C�   >\)   B�  >��>p��B(��@�  D�` A33?Vȴ   >��m>ٙ�?rn�?!%         @�        A�  ?�   =o>o��D��          >M��@�     A�  B�  A(z�@�  >Ƨ�F��UB�G�B�     ?L1B�     @��?�{@�C�G��ÿ��Ef}ţ+�G?}FP�iF��*ƀ�nE^���ƫ�]G?��G-��G�b7F
�QƯ3G��DK�|��}�A��ňV�	��F�VD5�$C}��ݦ�ŀo3��¼�"FG$եƵ9qD{UX�{������D?�5F�@��@a)�B�GG�)�/�������ǘ%ƅY�f�Ƹ$��=�CȰoF��F�quE�� �	�wF�&*Ʀد�Tp�G0O���pD=qF�19ř��F���Ųj�F�hL       split_indices[$l#L       }   
            	                                                              	               
                                                     	                     	                                                                                                                                                                                                                                                                                        L       
split_type[$U#L       }                                                                                                             L       sum_hessian[$d#L       }F�` Ey� FNL E� D� F Ep� D�� D@ D� D�� Fd B�  E!� D�  D�� C�� D@ B  C�� CW  D`  C�  F� Cy  Bt  B8  E  C  Ch  D�  Bl  D�� C�� BP  C�� B�  A@  A�  Cr  Bt  B�  C  DD  B�  B(  C�  F� C�  Cq  A   A�  B0  @@  B,  D�  D�  C  A�  A�  CW  C@  DR@ A�  A�  De@ C  B�  C>  A  B,  C�� C  B�  @�  A  @@  A`  A   @�  Cl  A�  B   Bt  @@  B�  BP  C�� Cʀ B�  B<  A@  A�  A�  C�  E� E�` C�� B�  Cf  A0  @�  @   A0  @�  A�  A�  A�  A`  D�@ A�  Ce  Dj� C  A  AP  @�  AP  @�  CP  @�  B�  B�  DP� @�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       125L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       iBL�F ��ğ�xG�b�E�O���yCDE�bF��EH] �J��F:�K���VƠ��TL`Eq�Ə\�F�TjG��kF"s�Ez�n�GZ�EC �F�~+E�3Ơ5pǑ�J�@"���[�%��; E�lmDQOU�IW�=�\F=/!F��L�]��ŏ�7F�4�FS.�GY�r���F���ƷZ�GP�0ƿN1Ǽe�G�ƍF�GdsC�n����8Ƹk�Ƿv��$v�F(���>2D� ā�E�ll���tE��ŕl���CD5������FզmE���G:�oE�;��1�,��i�F�����e�EF���f	F&P�D���C�]�G���F6H�N,��=�����F���EQV�ź�8GA��G�6�F)-E���e!Fm}��M��� �IGi�Gťz��3�8�8��@~/FIy�D�a��{6�E]�]L       
categories[$l#L       =                                   	   
                      	               
                      
                                     	   
                                     	   
            L       categories_nodes[$l#L                    	               !   &   1   7L       categories_segments[$L#L                                                                              !       "       0L       categories_sizes[$L#L                                                                                           L       default_left[$U#L       i                                                                                    L       idiL       left_children[$l#L       i               	                                 ������������   !   #   %   '   )   +   -   /   1   3   5   7   9����   ;   =����   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c   e   g������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       iR.�KRj�R A�Q��JQ��xR�u�RsglP��NP�upQ.8�Q���R�R�S#R='�Ro��N��Y            Q<T�Q*��Q��RH�jR�DR#�\R+I�R��Q���R��~R/FRl�:Lz�>    Q��Q+��    Q9G�Q��]R �pR�R�Z�R�*ER�x�R�ZR�i�QzS�R!��RMeR�=�R8�Qy9R�~�RۨQ���Q��S��Q�m2                                                                                                                                                                                                L       parents[$l#L       i���                                                           	   	   
   
                                                                                                               !   !   "   "   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8L       right_children[$l#L       i               
                                  ������������   "   $   &   (   *   ,   .   0   2   4   6   8   :����   <   >����   @   B   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d   f   h������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       i   <�   >hsB5\)@���>���Bb�\      AP     ?3��B�33      F�TjG��kF"s�B��D� ?�%>��R>9X@{�B9��>&�y=��`=��mD�� ?��T   �IW   B.��F��LD�` A0     ?���=�`BB  B<  B;�\B�  @���A�  >��jAp     =P�`>�-A�  B|ffA0     @�  D� ā�E�ll���tE��ŕl���CD5������FզmE���G:�oE�;��1�,��i�F�����e�EF���f	F&P�D���C�]�G���F6H�N,��=�����F���EQV�ź�8GA��G�6�F)-E���e!Fm}��M��� �IGi�Gťz��3�8�8��@~/FIy�D�a��{6�E]�]L       split_indices[$l#L       i      	                                                                  
               	   
         
                                                       
                                                                                                                                                                                                                             L       
split_type[$U#L       i                                                                                             L       sum_hessian[$d#L       iF�` E  Fg@ A0  EP Ey  F(� @�  @�  D)  D�  E) D�  D�` FL @�  @   @�  ?�  C�  C�  DT� DW� D� DG  C)  D�  Dh@ CJ  E�� E�� @   @   C   C�  @@  C�� D� C�  D3@ C  Dl  Dq@ D?� A�  BP  B�  B�  Dz� A�  Da  B  C&  A�  E� E�� Dy  ?�  ?�  A�  B�  CQ  B<  C2  B�  D� A@  C~  @�  C�  CY  B   B�  C�� C� C�� D#  Cn  D  A�  @�  A@  B   B  B�  B   B�  Dx� A  @@  A�  B�  DL� A   A�  C$  @   A   A  E� B�  C�  Ea� D9� C}  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       105L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       _BfrZ�@ۉDW����w���DD:YG���C4 �
����]�yt�D����uwRG�%s�坑G!���i�D��^�ǀ��$Ek�\�Ɖ��G:çĩ��E�RǠ�/m(G��EGyGvp<�fug����G�*F� u����+#���RoET2?�{���UM�ޗ�G������CS�5Ƈ��Eou/G���å�9��Jn�G��|G���gE�?�F��g��M�z��F_�D�*4D���F)���SRƢe�ŅL�Ɩ��&*��/mECbb�(R��x?����9�nF��2��DyM�G ��D�e4�A����6gD����ة�E��]���E���C��^F�'\E����
�|��Y��x�Q<�E06����*F�uE`@�L       
categories[$l#L       '                                                 
                            	   
                           
               L       categories_nodes[$l#L       
                  %   +   -   /   0L       categories_segments[$L#L       
                                                         $       %       &L       categories_sizes[$L#L       
                                                 	                     L       default_left[$U#L       _                                                                                L       idiL       left_children[$l#L       _               	                           ����         !   #   %����   '   )   +   -   /   1   3����   5����   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [����   ]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       _R�(Q)�R�QB�Q&�Q�^�Q�)�P�w�P���Q4� QI�R+U@R��QP�<    PJ[�P���P�h0P��P�k�    Q1YHQ&�oRhJ�R��Q�@XR>,CP^1�    P��    PD�NP�N�P���P�O@��P�7�P�CP��P̡(Ph��N�A�R<MR���R_�&RĪP�l�P5�@Q�A�    Pd�                                                                                                                                                                            L       parents[$l#L       _���                                                           	   	   
   
                                                                                                                 !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   3   3L       right_children[$l#L       _               
                           ����          "   $   &����   (   *   ,   .   0   2   4����   6����   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X   Z   \����   ^����������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       _@   >,1A�  D�@    D�  @n�R   >J��C  B  D�� >��B�33�坑?ƨD� =t�   ?��9�\�D�  ?>5?   B���B�=qA   D�� Gy=m�h�fug   B   >\(�BH  >q��Bff   ?���A�  @CoD�  @�   @=p�   D��       >�/G��|By33�gE�?�F��g��M�z��F_�D�*4D���F)���SRƢe�ŅL�Ɩ��&*��/mECbb�(R��x?����9�nF��2��DyM�G ��D�e4�A����6gD����ة�E��]���E���C��^F�'\E����
�|��Y��x�Q<�E06����*F�uE`@�L       split_indices[$l#L       _                                         
          
            
          
                                    	      	          
                                  	                                                                                                                                                                                   L       
split_type[$U#L       _                                                                                     L       sum_hessian[$d#L       _F�` D�  F|` C  D^� F| A�  B  B�  C�� C�  Ft� C� A�  @   A   A�  B�  A�  C�� @   C�  A@  F, E�� A�  C�  A�  @@  @�  @@  A�  @�  A   B�  A�  A   C�  B�  C�� C]  A   @�  FX D]@ E�X C�  A�  A0  C�  @   A�  @   @@  @�  A�  A  @@  ?�  @�  @   B�  A   A   A   @�  ?�  CB  B�  A�  B|  C�� @�  CE  A�  @�  @   @@  ?�  E�0 EY  Ci  D#  DB� E�  B�  C�  Ap  @@  @   A  C  C�  AP  @@  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       95L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       }B�H�.�lE&��E��{�s�}�m�E�E�F���	@����~�w�2S��F
�]��G:9E��l�IYaGНg�u/ō�X�,YF��p��pE�>�G�w�wG<ͻE������iǢ�GV�E=[H f�}iqH:YH4U�F���ƍ�%G�b�/!�}k��4W:G��-G+�@E�RHFO��ǉKF��m�7H/ƴ��� ��Gs�aF���G���FѤƅ�E�������YF�j���7�k�FsHF��.�0�UFZK]GJR�FN���'����(GpT8�1gGm�kF�hŴ�Fm1�Ŝv;�I	F��D�U��;���mE���ļ���d��FaiGY�\Ɛ�EH4F���0]l����
U�E��GS]Xǆ|�Č#�F�`�G�Ny�|:�E�C�Ʋ�����P9GF��Ʊu|F����BaG2���v�gE��cF5���~�d�FFw{�߄i�\�>�l|�/Ʃ�Fx�jL       
categories[$l#L       B                     	   
                               	   
                              	                                      	   
                                           
                                  L       categories_nodes[$l#L                         "   #   $   %   &   )   +   7   8L       categories_segments[$L#L                      	                                    .       /       <       =       >       ?       @       AL       categories_sizes[$L#L              	                                                                                           L       default_left[$U#L       }                                                                                                      L       idiL       left_children[$l#L       }               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W����   Y   [   ]   _   a   c   e   g   i   k   m   o   q   s   u   w   y   {��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       }QQ�{�R&�0Q�u�Qw��RE�RO�PR/WPR �}Q�N�RSR�R'�R��RRG]R��Q�cHQ�SXQ_.�Q���Q��vQ�X�Q��R��R�fQ��:Ri�R�;fRhY�R#inR@�=P� �Q�},Q��>N�0 R�^QR��NS O��R��Q {WP�m�Q\�Q�3    R �]Qk�5R'm�RpR[=@R�EQn|P2r�Q�W Q̤�R
fFR�m8R~"�R�tRy-Q��4RE��Q���                                                                                                                                                                                                                                                        L       parents[$l#L       }���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <   =   =   >   >L       right_children[$l#L       }               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X����   Z   \   ^   `   b   d   f   h   j   l   n   p   r   t   v   x   z   |��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       }BP  ?z�H>���?��>���@�        ?�=�"�A�  =��=ě�=�P@�  @@  ?�PBNG�??$Z@@  A�  D�     @XQ�   A�  B�B�   @Ϯ?I�@   B#
=BF��               ?;d>;dZ   =ě�   G��-BI��=ě�>��>��m@R�\@_\)>�r�D�@ >D��>��      @�  >�X?2n�B{��>�?�  ���7�k�FsHF��.�0�UFZK]GJR�FN���'����(GpT8�1gGm�kF�hŴ�Fm1�Ŝv;�I	F��D�U��;���mE���ļ���d��FaiGY�\Ɛ�EH4F���0]l����
U�E��GS]Xǆ|�Č#�F�`�G�Ny�|:�E�C�Ʋ�����P9GF��Ʊu|F����BaG2���v�gE��cF5���~�d�FFw{�߄i�\�>�l|�/Ʃ�Fx�jL       split_indices[$l#L       }               	              	            
                  	                                      	                                 	                   
      
                                       	                                                                                                                                                                                                                                                           L       
split_type[$U#L       }                                                                                                               L       sum_hessian[$d#L       }F�` F\ Fd D>� E�� D�` E�p C�  C�  Ec� Er  Db� C�� E�H EBP C  C�  C�� A  DF� E2  E_� C�� C/  D6� Ap  C�  CE  E�  E7� C(  @�  C  C�� @@  C�  @�  @�  @�  D=� B  A�  E0� E_� ?�  B�  C:  B�  B�  C�  C�� A   @�  C�� Ap  C  B@  Ey� C E(� Cs  C  B  @�  @@  B�  Bt  C�� B  @   ?�  Ct  A�  @@  @   @@  ?�  @   @@  D<@ @�  Ap  A�  Ap  @�  B�  E)  DD@ E.� B�  @�  A@  C.  A�  B�  B8  B  C�  A   A  C�  @�  @@  @�  @@  B�  CW  A   @�  AP  C  @�  B,  D�� E0 B4  C�  E� C  B�  B�  B�  A�  @�  A�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       125L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       uB)6�E,��F|�E���ñ���˜�EL�F���D
���+V�G����o�F5a�6ӡF^��F�� ��9D�Hs�h�nD�&�(eGu��G%�Y��džEG��Ō�uF":�� g�H��F9���щNF�b���?��*[�Å��G���"+��aDΰ�H��G"���Zv���G����dm��Qӣ���d2$F|P�G����ss��u�O��Ghv~FzƗ����Hp2�F�м����Q����4E��)FK���I�Gn��py:F_ʴD�[�3�F�&}E��@�G^bG �ǂ=��R�D/W��_GT?���ZF�V�ƫ��Ƈ���5KG>dE�ZMš��F�cA��;��%À_R�9d� [���P�E�� Ǫ7\Fj��G<&Zœ��F��E?�]�$�-FHG�JxC�oF� sħ� �3�Ʒ���dw�G��Ff@�F5�D*�E�ƨ6L       
categories[$l#L       7                                 
                                  	   
                        
                  
                                              	   
         L       categories_nodes[$l#L       
             	            .   0   :L       categories_segments[$L#L       
                                                         &       *       +L       categories_sizes[$L#L       
                                                                      L       default_left[$U#L       u                                                                                                   L       idiL       left_children[$l#L       u               	                                    !   #   %   '   )����   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S����   U   W   Y   [   ]   _   a   c����   e   g   i   k   m   o   q   s��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       uQ�~}R��Q��R�ЛRB��RY�R�:R�|�R>7R#��Q��R
��R� R2��R{�RH[�R�8�R	�RݪR�/RX��    Q��nR��Qˤ�Rw�RG�R�P�RV�:RTؒRO(Q���R?jlR]hQ�_�Q���R0�Q��Q��lRK�>Q90�R_"�Rf2    Q���Q��dR�RU�R>�R1��Q�~lQ�     RP�dR���R1�Rb*�O��Q�k�RO�(R"
H                                                                                                                                                                                                                                L       parents[$l#L       u���                                                           	   	   
   
                                                                                                                                   !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <L       right_children[$l#L       u               
                                     "   $   &   (   *����   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T����   V   X   Z   \   ^   `   b   d����   f   h   j   l   n   p   r   t��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       u   @B�\      CW
B�  ?"JA0  B�     @���=�7L   >J=�P=#�
@�  B�  >�B`  D�� Gu��D�  B���   ?��D�` =�"�   >oD�� @�  Bp  ?>��?��B�  A   >���D�� BD  @�  @P��=�Q����D�  A�     A"{   @�  >��?�/�u�O?�B��{?�/@@  =��#   ?L1@o�Q����4E��)FK���I�Gn��py:F_ʴD�[�3�F�&}E��@�G^bG �ǂ=��R�D/W��_GT?���ZF�V�ƫ��Ƈ���5KG>dE�ZMš��F�cA��;��%À_R�9d� [���P�E�� Ǫ7\Fj��G<&Zœ��F��E?�]�$�-FHG�JxC�oF� sħ� �3�Ʒ���dw�G��Ff@�F5�D*�E�ƨ6L       split_indices[$l#L       u                                                  	                                                                     	                                            
                   
       
                                                                                                                                                                                                                                   L       
split_type[$U#L       u                                                                                                           L       sum_hessian[$d#L       uF�` F� E�  EE@ E�� E�� E,� D�  D�` E�  A�  Ev` C�  D�  DH� D�� B�  D�` B   E�� D�� @�  A�  C� EYP C  Cu  D.@ D�  A@  DE� A0  D�` B�  A�  D�@ B�  A�  A`  E�� @�  B�  D�� @   A�  C�� B�  E� D�� B�  B0  Cq  @�  D  C	  Cǀ DX@ @�  A   D*  B�  @�  @�  D� C� B�  @�  Ap  @   D�  B�  A�  B�  A�  @�  A   @�  E�@ A�  @�  ?�  B�  A`  B�  D�` @�  A0  C�  A  B�  BD  E� B�  C�  D;� B�  ?�  A�  A`  C$  B�  C΀ C  B�  A0  C�  Bl  C�  C�� ?�  @@  @�  @   C�  C�  Bp  BL  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       117L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       gB�E��EĂ�NG�i�E���D�8��@�Fcy`H)ӀƭE��k�Ɏ\E�YED����,mHƔ)lG-��Gf�F��A�w�JQE�F�_CL^��e���X�qF3xk��vG���ɠ��������:{FsF`EN�'��F���ƍ�7Ǧ�CG�l�E�3�Ǣ�GF���ű+E}��G��l�{2�F�5�ۣ�E�GF��$C%�y�@&G�3��*Y��l�F ��G�O����E�����rWF�IK�	�'GIhcE���F�nDH@�f ��o'�F!�����oC�KGńD٤�łGUYġ��4�����FN�s�.��D��Cb?�E�. E�T>F���큈EU
��/���QZGAˀFn��ƒ`�FKRa�@��V��F�JŪw���?GrP��_�Gc|
L       
categories[$l#L       F                       	                                  	   
                                           	                                      	   
                                             	   
                        
   L       categories_nodes[$l#L                                $   (   )   -   .L       categories_segments[$L#L                             	                     $       %       &       2       3       4       AL       categories_sizes[$L#L                                                                                           L       default_left[$U#L       g                                                                                   L       idiL       left_children[$l#L       g               	                                    !��������   #   %   '   )   +   -   /   1   3   5   7   9����������������   ;   =��������   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c   e��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       gQ��Q���Q�*fQ�!�Q�1�R!|PQ�7|O�ZPU�pR' Q�yiR@�RI�?Ro~�R��M�&XM��        Q�#�Q��Q�
�R) lR ��RF�RR��R@�`R zaQ���RTYR���                R	��Q_5�        P�*�Q��jQA�JRWQR$ɿR#�Q��Q�2�Q�K�Q��hR'Rb��Q��LP��QR�@P�RbR�R���R:o�R1�,                                                                                                                                                                                L       parents[$l#L       g���                                                           	   	   
   
                                                                                                               #   #   $   $   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   :   :L       right_children[$l#L       g               
                                     "��������   $   &   (   *   ,   .   0   2   4   6   8   :����������������   <   >��������   @   B   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d   f��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       g   <�A   >hs=��
@�     @@     @�  B�  @�  @�  AP  B�        Gf�F�      =�{=�1?9X>�ffD�@ >�9XB�  @�  D�@ =�h�����:{FsF`EN�'>��m   ƍ�7Ǧ�C@�        A$��>�K�?��      >��F@��B  B�k�@�  B�R?hsB���B�  ?�n�=���C  E�����rWF�IK�	�'GIhcE���F�nDH@�f ��o'�F!�����oC�KGńD٤�łGUYġ��4�����FN�s�.��D��Cb?�E�. E�T>F���큈EU
��/���QZGAˀFn��ƒ`�FKRa�@��V��F�JŪw���?GrP��_�Gc|
L       split_indices[$l#L       g      	                                                                     	   
                                        
                           
                 
                                                                                                                                                                                                              L       
split_type[$U#L       g                                                                                           L       sum_hessian[$d#L       gF�` E  Fg@ A0  EP F0� EZ� @�  @�  B�  E F� E$0 D�� E� @@  @@  @�  ?�  B�  @�  D�  C�  E� D�  C�  Ep D�  A�  E� BP  ?�  @   @   ?�  BP  B0  @   @   @�  D�@ A`  C�  E<� E�� A`  D�` B�  C�  D�� C�  D�� @�  A�  @�  D�  C�� A`  B  A�  A�  A  B  @�  @@  B�  D� A@  @   C�  A@  D΀ D�� E� Cˀ @�  A   D,� C�  A�  B�  Ce  B|  D�  CÀ CĀ B�  DQ� C�  ?�  @�  AP  A   @@  @@  D�@ C^  C~  CC  A   @�  B  ?�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       103L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       oAފ�ě��Eyt��N`��+#���X�E��D1��̕��ԥ?ǝU�Ʈm����G�Z�E����"��Fh���1��E�	�� ��4�"�ͬ���u�G�(����+�aU>�`�)G$2�H��~E6i�G+M�ņ�*EgzB��G/k������
>Z���FY��揟F��F���H��ǀ����G_� ǌlG8�J�	��G������E�[ZǈPG�^��5�ōO�H�!�Fu��Ca�G�I��	K��w���I7F�'DMӧD��b�;�E�2QF�o��#�Eݰ�ŭ��Ʋ;ƙ���2��D�-eF���E�B-�|�eFVl����ƅ$kE�ؔ�$���QMƓ-��E�|F�j}E���=;�����GAD�E:F3_��2HXD^�gƹ��G�ibF)����p�F��-Gˆ
ċ#�F/'���6Dǲ�G�Ą!����C�lL       
categories[$l#L       >                                                 	   
                                            	   
                                           	   
                                    	          L       categories_nodes[$l#L             	          ,   -   .   1   2   6   9L       categories_segments[$L#L                                                         #       $       1       8       =L       categories_sizes[$L#L                                                                                    L       default_left[$U#L       o                                                                                              L       idiL       left_children[$l#L       o               	                                    !   #   %   '   )   +   -   /   1   3����   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O����   Q   S   U   W   Y��������   [   ]����   _   a   c����   e   g   i   k   m��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       oQ���RXl�R��Q�%Q�$�Q��QR�0`Q��RZ�Q(4Q��Qq(QvDR�[R:	^R=R��*RE�R�pP�P�A�P� Q:6�P��RQ��P0��    R��Q�8Q���R� R'�R�*�Q���R��9Q�ػRB�XQ���R&�pP��PH_�    P�ĘPH��P�%`N�w�O3�        P���QB�n    O���Q��vQ(��    P�@R���Q���R���Q���                                                                                                                                                                                                        L       parents[$l#L       o���                                                           	   	   
   
                                                                                                                                   !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   *   *   +   +   ,   ,   -   -   .   .   1   1   2   2   4   4   5   5   6   6   8   8   9   9   :   :   ;   ;   <   <L       right_children[$l#L       o               
                                     "   $   &   (   *   ,   .   0   2   4����   6   8   :   <   >   @   B   D   F   H   J   L   N   P����   R   T   V   X   Z��������   \   ^����   `   b   d����   f   h   j   l   n��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       o?"J?L1D�� >� �B�G�   D�@ A33@�   A	��=���B�  A   B�  >9XA�  B�ff=���D�  B  D�� @~�+   =��wB��`�)?+C�A�D�  ?���?�   A$��>���?.�@�33@@  B���B@Q�@kC�F��Bz=q@�           G8�J�	��      E�[Z>hsB�     ōO�@@     ? �@ǮD�� �w���I7F�'DMӧD��b�;�E�2QF�o��#�Eݰ�ŭ��Ʋ;ƙ���2��D�-eF���E�B-�|�eFVl����ƅ$kE�ؔ�$���QMƓ-��E�|F�j}E���=;�����GAD�E:F3_��2HXD^�gƹ��G�ibF)����p�F��-Gˆ
ċ#�F/'���6Dǲ�G�Ą!����C�lL       split_indices[$l#L       o                                                                                                                                
                                            	                    	                                                                                                                                                                                                              L       
split_type[$U#L       o                                                                                                    L       sum_hessian[$d#L       oF�` FKp E�� FIx B�  C	  E|� F� E*� B�  B  B�  A@  B0  Ey� F� D@ D�  DJ@ B  BL  A�  A   @@  B�  A  @@  B  A   ErP B�  E�H E�� C�  C�� Dɠ C�� B�  D0� Ap  A�  @   BD  Ap  AP  @�  @�  @   ?�  @�  B�  ?�  A   A�  AP  ?�  @�  D(@ EH@ B�  B  E�� B�  B�  E�� C^  B�  C;  B�  D�� B�  CZ  B�  B  B�  D$� B@  @�  A   A�  @�  B8  @@  A  @�  @�  A  @�  ?�  ?�  @�  @@  @@  A  B�  ?�  @�  A�  @@  @�  A  ?�  @�  C�� C�  D�� D�� BT  B  AP  A�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       111L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       {A�˗�	%OD�EE��<�/�BD�?����FG,z��ٔ�Ś-ƋdB�8zF	��G���"�{G�XKŘ�9�@h�F�3����p�SH�.�&��dFyā�+3�F��v�1vyFvO�Ho xGkƺ�I��G'�G,n�F�z=��D0���E���G��sE!=��Y��`�š�cFt9���C^ŃtHFId���E�0�G���DP�:�	OF��ǻ�lF����b7Ǌ�oGN�IH���FP����R�HEE��9��oEL<F�LY�+�zE�:��é�gE�W�_�E�O�Ű*�Gm�E&\�F3��Ň�EPD:���ą�MƟt�D����VZ�F��vċ�D��*����B�6��c��F/rJ�1��ď��F�R�B+E�G(���)<��5�E��>DcP���NGE�!�F�2Ɔ������<G8�I���%���F���$*E�t�G|�FӫLG��F�����Ex��G�������֢;�'�F�L       
categories[$l#L       C               
                             	   
                                  	   
                                                           
                                  	   
                            L       categories_nodes[$l#L       
      
         "   #   %   0   7   ;L       categories_segments[$L#L       
                                                   %       1       =       BL       categories_sizes[$L#L       
                     	                                                 L       default_left[$U#L       {                                                                                                          L       idiL       left_children[$l#L       {               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?����   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c   e   g   i   k   m   o   q����   s   u   w   y������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       {Q���QΠQ���Q �_P��lRE�R+:P��P��P�U�P�� Q��ER���R�W�RAP�� O���P�-�Q$Pw0<PN�P�?/P��|RS�R�tR�<�Q��R�Q�dR��GRH�oOݤ4    N���N%żP�q�P�4OԬ�P}�PO}��O�P��P� P(�,P�P�P�`P���R��R���R84R�RRs�8RqF�RM��QxaBR>��R��N�B     Q�T�Q�cRS `R E
                                                                                                                                                                                                                                                L       parents[$l#L       {���                                                           	   	   
   
                                                                                                                                 !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   ;   ;   <   <   =   =   >   >L       right_children[$l#L       {               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @����   B   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d   f   h   j   l   n   p   r����   t   v   x   z������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       {B   D� D�� >�A�   D�  ?��R>��>x��>_;d   =��`   ??}=��>vȴ@�  >��=Ƨ�>R�?+�>�o>	7LB��{B�\B�  ?�  @      Bfff>���?�  G,n�A�      ?!%   >���D�� @   ?^�RD�  =���=�{A�@,�>��   B�  ?�G�A�  ?�G�B�  >�o   >��DB�
FP��   >���=�"�@�  EL<F�LY�+�zE�:��é�gE�W�_�E�O�Ű*�Gm�E&\�F3��Ň�EPD:���ą�MƟt�D����VZ�F��vċ�D��*����B�6��c��F/rJ�1��ď��F�R�B+E�G(���)<��5�E��>DcP���NGE�!�F�2Ɔ������<G8�I���%���F���$*E�t�G|�FӫLG��F�����Ex��G�������֢;�'�F�L       split_indices[$l#L       {                                     
          	         
      	         
                                             
                      	                                         	                                                                                                                                                                                                                                                                   L       
split_type[$U#L       {                                                                                                                 L       sum_hessian[$d#L       {F�` Dl� F}� B�  DN� Fj D�� A�  B�  CӀ Cɀ FF� E B�  D�� A�  A   B�  A�  A�  CȀ C{  C  C�� F@� D�` D� B�  @�  B  D�� A`  @@  @�  @�  A�  B  @�  A�  A0  A0  C�� B  B�  C,  Ap  C	  C�  B4  F"l D� D�� A�  BD  D@ A�  B�  @�  @   A�  A@  C�  DF  @�  A   ?�  @@  @@  ?�  @�  A�  A�  A�  @�  ?�  A   A�  @�  @�  @   A  C  CY  A  A�  A   B�  A�  C  @�  A0  B�  A�  A�  C�  A�  A`  F� C�� D�  Dc  D�  C.  A�  @@  B   A  C�  CW  A0  A�  B   A�  ?�  @�  @�  A�  @@  A  BL  C�� D,@ B�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       123L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       KA�8C%f� W��RE�E�����>Ƨ���C�O�E�@}H kQ�p����SƁ�x�=zJ�S�-ƻ�~��x�F-1XFW�Ť��H�Bl����K�F/G�E��F�a������G���D;
��.�F�(����G^E���<
�F�>�GFa�FW�TE�����!Ű�ǂ�
����F��GguD���Ę|�D�Ɨ�~ū��G%^F-����5E�89�T��Fzs;FA4l�������Fe�Gf�E���D<��FC��E�'�ŢdrF:�fņ��E�ŧ/����fŰ�Ɓ��E�%�L       
categories[$l#L       2                	   
                               	   
             
                               	   
                                           	   
         L       categories_nodes[$l#L                
               !L       categories_segments[$L#L                                                                $L       categories_sizes[$L#L                                                               L       default_left[$U#L       K                                                               L       idiL       left_children[$l#L       K               	                  ��������   ����               !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C����������������   E   G   I����������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       KQ��Q�c�Qs�Q�m�R"�DN� Q7tR� Q�؄Q��.QB,        P�b�    Q�P�Qɖ�Q�cR?v�RA��Q��QN}� N�;.Q	�Q~�Q�NRcoQ��4M:� R
��R��lRkK�RLcS8R �Q�[QХ�                P�P��(P��                                                                                                                            L       parents[$l#L       K���                                                           	   	   
   
                                                                                                                       !   !   "   "   #   #   $   $   )   )   *   *   +   +L       right_children[$l#L       K               
                  ��������   ����                "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D����������������   F   H   J����������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       K@��;?�>�\)@�  A�     B�     A33@���   �p����SB�B��=zJD�` A�     A�@@  @c"�A�     @\�@�  =�t�B�G�      >�/E}  @�  A�     @�
=??}?��GFa�FW�TE�����!>�bN@   @�hF��GguD���Ę|�D�Ɨ�~ū��G%^F-����5E�89�T��Fzs;FA4l�������Fe�Gf�E���D<��FC��E�'�ŢdrF:�fņ��E�ŧ/����fŰ�Ɓ��E�%�L       split_indices[$l#L       K   
                                                                 
                	                                                                                                                                                                                        L       
split_type[$U#L       K                                                                   L       sum_hessian[$d#L       KF�` F�� B�  Fbl E%  @�  Bx  D� FF< E$` A   @   @�  Bt  ?�  D�� C� F9( DQ@ D�@ DC  A   @   B   A�  D>@ D  C� @�  F� D�  C�  C�� C�  D�@ D@ C#  @�  ?�  ?�  ?�  A�  A�  A�  @@  @�  D=  C�  C  B�  C�  @@  ?�  F\ C�  D�@ B�  C�  C*  Cw  B�  A�  C�  D�� B�  B�  D  B�  Bl  @�  A�  A   @�  @�  A@  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       75L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       kA�~E_RAĤKKǸ��Er��Ç�K��|�
��	�3ZE�-jħ&�F�n��-|č��F=�EƓ�}�9�|�U�TF%	�ٽ�Ez,�F��T�G�4+wE��GE���TYF/U
�q�Ez5�ĭ�����Ej'hHk�ķ���e�>E�wYŬ��GL�HE8;�ϭ�GD��o8HG�Fܬ�ƍ\G�&�F{��F���ǉ�G�"��l�?�G�~ǃ�E��� [M�� F/M;�9���'GQ��^�G%d��:c���(TD���FSg�E h��aKG!]�F	��E�qS�}��E`�éS�EyrG.��t"���zZEG�F�χE�D�F��FF��� ��FڠG?E�F��X��W�͋sFMƆ���2wE��GX�GZ�Ƌ�BNϖơ�xG��V�7Θ��`F���E�xz��3L       
categories[$l#L       F                                                           
                  	   
                               	   
                                                                                            	   
         L       categories_nodes[$l#L                                   '   +   /   0   2   5   6L       categories_segments[$L#L                                                                              (       -       .       2       4       :L       categories_sizes[$L#L                                                                                                                L       default_left[$U#L       k                                                                                      L       idiL       left_children[$l#L       k               	                              ����   ��������   !   #   %   '   )   +   -   /   1   3   5   7   9����   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c   e   g   i��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       kQ��.R�Q�y�Qk��Q��5RRvR�%�O�'yPzR%�R��Q���RU��RXy�R^e    N_�h        R��R[ڦR�lR1X�Q�SR7��RF�ER�G�R���R�IR�O
RJH�à    Q��ZQ�mR
�Q�r(Rw"Q�=�R�5�RM�Q��~Q�8Q�a�Q.H�R�RјRnnDRu�;R�OR8R>TR7"�R�*Ry`�RF�%R:�                                                                                                                                                                                                        L       parents[$l#L       k���                                                           	   	   
   
                                                                                                               !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8L       right_children[$l#L       k               
                              ����    ��������   "   $   &   (   *   ,   .   0   2   4   6   8   :����   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d   f   h   j��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       k   D�` B�\>��^>��hB�  >V      >]/B     @��>��^B�  F=�E   �9�|�U�T@�        @�  C  E}     >��=�h>��Bd  >�Q�Bff���>&�y>I�^@�  B�ff@c"�?|�   B�  =�C�>���   >���D�� >o      B�     D�@ =� �      @�  @@  � [M�� F/M;�9���'GQ��^�G%d��:c���(TD���FSg�E h��aKG!]�F	��E�qS�}��E`�éS�EyrG.��t"���zZEG�F�χE�D�F��FF��� ��FڠG?E�F��X��W�͋sFMƆ���2wE��GX�GZ�Ƌ�BNϖơ�xG��V�7Θ��`F���E�xz��3L       split_indices[$l#L       k                               	                                                             	   
                            
                       	      	                                                                                                                                                                                                                                          L       
split_type[$U#L       k                                                                                            L       sum_hessian[$d#L       kF�` E�� FB� A`  E�@ F)� D�@ @�  A  D � E�0 F � D@ C�  D�@ ?�  @�  @�  @   Cb  C�  Es  C�  F� D� Cƀ C$  Cj  B�  C&  D�� @   @   CY  A  C  C  E*0 D�� C  C  FT B  Dn  B�  CP  C=  Bp  B�  B$  CA  A�  B@  C  A0  A�  D�� ?�  ?�  Bx  C  @   @�  C  @�  B�  B  E$  B�  C�� DG� B   B�  B�  B  C�� Fx A�  A  C� C�� B   B  C(  B   A�  C+  A�  B  BL  BT  A  B   C(  A�  A   A@  @�  B,  B4  B�  @�  @�  A�  A  D� C�� L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       107L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       uB]��6�D�D_�Yz�G��F�>Co3��E�Rǫ#F/ˍG��Gg-Đ3sD��!�~t!��IfD��
ƚ���DT�GXG��
6�H{�NGM�F��EG�}���%F�1�D�F��?GF�Ƨ�>Ɗ0�BئF��?�`>OGX�#�hPǮ u��� G���ƅ�0�WB2Ff��G�1�Ft�G�k��8�`E���GTGzS�Heh�Ŋ���+z}Gw��B��L�D�WG�
F=A�F���G�-F�`��ǈ��ļ�K�@��,s�EF<FcS4D��D���ő��F�4�D�B��zL���aF�EŐ6��#�ƞ��Œ� FBJ�G_��F!�E�*�$���p�E�:Fْ���F���ťunG��[E���F�}��A����qE��+G?�
DN�GƝ�{ņ��F��lF8��C��PG9�ƽz�F
���s�TF�9Ċ��G)��Ec�W��\JF3���� %G�ݟL       
categories[$l#L       J                  	   
                                               	   
                           	   
                     	                                     	   
                                                 	   
            L       categories_nodes[$l#L                      !   "   #   $   '   .   <L       categories_segments[$L#L                                                  $       *       7       9       ;       >L       categories_sizes[$L#L                                          
                                          L       default_left[$U#L       u                                                                                                      L       idiL       left_children[$l#L       u               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I��������   K����   M   O��������   Q   S   U   W   Y   [   ]   _   a   c   e   g   i   k   m   o   q   s������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       uQq#�Q��Q��Q�z�Q��_R�� RݼQ��Rc�Q�B�Q��6R�
�R#SRA(R89Q̒R~y+QEQ3QM��P�%�P�
�Q}�NR��R�
�Q���RT&eR��R��fQ?�$R'�}R?��Q�H6R2�(R2�rO�9�P��u        QX/z    P"�$O���        Qw�O��R.��Q���R��R�ܞR+҂Rc�R���Q8C�Q�dKR/ �R��@R.�BQ�Q~2Ryo�S
�                                                                                                                                                                                                                        L       parents[$l#L       u���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   $   $   '   '   )   )   *   *   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <   =   =   >   >L       right_children[$l#L       u               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J��������   L����   N   P��������   R   T   V   X   Z   \   ^   `   b   d   f   h   j   l   n   p   r   t������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       u?;dC  ?I7LB�  @�   A�  >�?}   >,1D�  A�  ??|�A�  =8Q�@�  >�n�>�w@�  =�S�>�X      @�  B�=qB��q>���>gl�D�  >��B��q>ؓuB$              Ǯ u���    ƅ�0@�  >C�G�1�Ft�@P     =�@��?8Q�@�  B��@9��B�ffB�  ?�=�P>�S�B�aH>1&�   @���?*=qļ�K�@��,s�EF<FcS4D��D���ő��F�4�D�B��zL���aF�EŐ6��#�ƞ��Œ� FBJ�G_��F!�E�*�$���p�E�:Fْ���F���ťunG��[E���F�}��A����qE��+G?�
DN�GƝ�{ņ��F��lF8��C��PG9�ƽz�F
���s�TF�9Ċ��G)��Ec�W��\JF3���� %G�ݟL       split_indices[$l#L       u                                	                     
   	                            
   
                                                                                                     
                                                                                                                                                                                                                                        L       
split_type[$U#L       u                                                                                                          L       sum_hessian[$d#L       uF�` E�p F< E�` B�  D�� F&L E�� A�  B,  A�  C�  Dy� Fl D  E(� E� A@  @�  A�  A�  @@  A�  C�� B�  DD@ CV  F@ CK  B   D  D.� D�@ C�� D�� @�  A   @   @�  A�  @@  Ap  @�  @   ?�  A0  A  Ch  Bd  B�  A`  D3� B�  B�  C  D;� F� B  C%  A�  A   C�  B�  C�  Cu  D�@ D:  C:  C?  D�` DH@ @   @   @�  @�  A`  @�  @@  A@  @@  @@  @�  @�  @�  @�  B8  C:  B$  A�  Bl  A�  A   @�  D,@ A�  B(  A�  Bx  A�  B�  A   D9� A   C  F� B   @�  C  B  AP  A�  @�  @@  C�� B�  B|  @@  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       117L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       ABCf�@�-�G�h�Í��F8^	G2մG �A��ƒc�Fj%����GxS�bZ ��(�GR�G0����UG��ı �d]�E�I�F�I��bWD���G�K���+H	�]F��Ǫ�-Ɗ/�G���n~ƲoG���F%��ş���@GǬM���8�ŭ��õ.D�!�G�IF.:N�D��GJ�UGU���D�[�F�=��4r�ԋ���q�G3�hF~� Şi'E���Ǆ#ś]6��G+�����E�D	�L       
categories[$l#L       %                      
                                   
                                     	   
                   L       categories_nodes[$l#L          	                     #L       categories_segments[$L#L                      	       
                     "       #       $L       categories_sizes[$L#L              	                     
                            L       default_left[$U#L       A                                                        L       idiL       left_children[$l#L       A               	����                  ����                  !   #   %��������   '   )   +   -   /   1   3   5   7   9   ;   =   ?��������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       AQb �QZ��P�|Q���R 
�    P
�qQ��R��R'�XQ��lM'[�    Q�<�R8^DRj�R;s�RoUR8�`N��PH��        R	�6Q�O�Re�R[�Q��P���RY�>Q�'�R�^R<̂Q��RL��Mc�                                                                                                                    L       parents[$l#L       A���                                                     	   	   
   
                                                                                                                       !   !   "   "   #   #L       right_children[$l#L       A               
����                  ����                   "   $   &��������   (   *   ,   .   0   2   4   6   8   :   <   >   @��������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       AA�  B�  AP  @�  A`  G2մ?��B�  D�`    >�   �bZ          >t�jB�  ?F�y      E�I�F�I�@�  BP  >��?��>7K�B�  >�B�  @&=u?�\)?�n�   ş���@GǬM���8�ŭ��õ.D�!�G�IF.:N�D��GJ�UGU���D�[�F�=��4r�ԋ���q�G3�hF~� Şi'E���Ǆ#ś]6��G+�����E�D	�L       split_indices[$l#L       A                                                              	                         
                        
                                                                                                                          L       
split_type[$U#L       A                                                         L       sum_hessian[$d#L       AF�` F�P A   F� C̀ @   @�  F�� C�  C�  A  @�  @   F�h B�  B`  C^  C^  C4  @�  @�  ?�  @@  E�@ F70 A�  B  A@  B0  BX  C(  CP  A`  C  A�  @@  @   @   @   E� D� E�X E� A   A�  B  @�  A   @   B  @�  A�  A�  C%  @@  C(  B   A   @�  C  A   Ap  AP  ?�  @   L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       65L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       }BZVEC�ĩ+4�i�E�aF~����D��ƖʸEU+�F�q�G�k��)ƤJF��>hF��%�ǚA>�]��F�4LE
��G'�_�%-�G��D���EP��3_L�/���u��F>����Ŗ˶F��VƄ�������h�Ƃ��{"�Hhb(Ǩ�F�ߩ���{E��E]g�G�&�ś5Ǐ>�G�Hc�ƃ��H�ጝFfI��[��G25���v�ǲ\>H����^xF�Q�ƖW�ŌRoE;��EjJ�	LF���E�&�F�i����3GI*�;)?F�k�H+qF-�{ƙ��6��m�qG��0F���FDLc�%�F�PRE(�o���Ƙ��C��#E���Fo���۩@Fp@�Gp��IWVFkٗ�'�pE%��s��F�ܽG��AF�\,�]�F{�YG�zF]�{�02��%X���7F�oƘ]bGW��bE���=��RGK��E֊4ġ2��I��E3xmFr��C�h��b�D���	O�EL���D��L       
categories[$l#L       :                                     
                                                    
                                              	   
                            	   
         L       categories_nodes[$l#L             
         #   &   (   )   8   =   >L       categories_segments[$L#L                                                                        "       %       0L       categories_sizes[$L#L                     
                                                               
L       default_left[$U#L       }                                                                                                             L       idiL       left_children[$l#L       }               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c   e   g   i   k����   m   o   q   s   u   w   y   {��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       }QU�kR'O�R#;Q�$�RN>R_�R3R��R!��Q��RhM�R�O�Q��eR~�Q̨�Q�<.R�RF��Rnf8R#�>Q��3R�[�Q/�kR�G$R��Q`UTQ��Q�Q�Q�/R�Q��XQ���R�fQ;�R!s�Q��pQ�R	�O䑀Q���RXw�R	��R*�R$�R�d�Q�bQp^�Q�;`Rf��R�`�RN��Q��Q��pQ� z    Q� �Q��dP3l(Q�BARܕQ�1,R5��Rt��                                                                                                                                                                                                                                                        L       parents[$l#L       }���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   7   7   8   8   9   9   :   :   ;   ;   <   <   =   =   >   >L       right_children[$l#L       }               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d   f   h   j   l����   n   p   r   t   v   x   z   |��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       }@B�\>)��D�� D�� ?�P@�\)>��
   >o>B�\   @   B�     >C�@@  B�aH   ?WK�<�t�D�` D�� ?q&�A�  B�  >,1@$��>��R=��`>���?b>1'=��<�t�=<j   D�� B�33   >=p�      By33>�JB���@�  ?�G�>�"�A�  @�(�>O�Bd  Bv{D�� G25�>��7   BVff@�  D�� BW��      EjJ�	LF���E�&�F�i����3GI*�;)?F�k�H+qF-�{ƙ��6��m�qG��0F���FDLc�%�F�PRE(�o���Ƙ��C��#E���Fo���۩@Fp@�Gp��IWVFkٗ�'�pE%��s��F�ܽG��AF�\,�]�F{�YG�zF]�{�02��%X���7F�oƘ]bGW��bE���=��RGK��E֊4ġ2��I��E3xmFr��C�h��b�D���	O�EL���D��L       split_indices[$l#L       }                            
                                                       
      
      	      	                      
                                                                                                                                                                                                                                                                                                                                   L       
split_type[$U#L       }                                                                                                                  L       sum_hessian[$d#L       }F�` E�P F* D�� E�� D� F!� D@ D� E�� C�� C�� CQ  C�� F� C�  B�  B0  D� C�  E�X Cw  C  C  C2  C  BX  C  C_  D:@ F( Cy  Ce  B�  A�  A�  A�  D  @@  AP  C�� D�� EY� B�  C  B�  A   B�  BP  C   A�  B,  B�  BP  @   B�  B  @�  C[  D� C  E�X E� C#  B�  A�  CL  @�  B�  @   Ap  ?�  A�  A@  AP  CԀ B�  @   ?�  @�  A  B�  C2  Dx� B(  E!� D`@ B  B�  B�  A�  B�  A0  @�  @�  A�  B�  A�  B   B�  B@  A   A   B  @�  B�  A�  BH  @   B�  A�  Ap  A�  @@  ?�  CX  @@  C�� B�  B�  Bh  D�  E�P D�  Dc� L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       125L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       mB/<C���ƒ�8AŞ8F��B�ou3�S��C����a�OG3����jǗ�aF���)��͑�D`��ũ�!G����aMH�f-F�n�FL������,�ǰ�aF3=�D�3ƉLJF�\�Ɛ���h�B4�F(xk�n�rƽ��EP9�G���̪Ǜp5G:N�H�C2���bGE�zEI�GS*�)\�F�A)F/��:$�T�K��8�żlǃ�����Gj�R��GF��Pĝr��/���d��E��E��fŮ����[	E� 8��g�F�'I���rF��F�hS��(IƉ=�š�v�M�F�2�G8XNH��ZH��/{@E�AF��Ex��t�F�$�Cc6g��8��UK�KE�G �nE�tDr�4�v��Ƈ���ehg�8��.��EQ����A�ͻz�w&5F'�F��E����]��[�O�`y�F7W$ǅ<�Ŵ�L       
categories[$l#L                                   	   
                                                                    L       categories_nodes[$l#L          	   
               $   '   (   1   4   5   6L       categories_segments[$L#L                                                                                                   L       categories_sizes[$L#L                                                                                                  L       default_left[$U#L       m                                                                                        L       idiL       left_children[$l#L       m               	                                    !   #   %   '   )   +   -   /   1��������   3   5   7   9   ;   =   ?   A   C   E   G����   I   K   M   O   Q   S   U   W   Y����   [   ]   _   a   c   e   g   i����   k��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       mQ�$ZQ��cQ%wzQo)�R�Q�XP�1QV�R\��S�Q^��Py!�M��P�C�Q��Q��Q���Q�K%R��REX�R>�P�ҔP�;ZN�E^P��        P��Q��QRB�P��$Q�^R�WQ��Q��Q�"DQ�
Qw6T    O��(P���Q}M�Q�7�P�;�P'� Q0w�Q�I�KK%     N`N�Y@P�˨OޞXP*��P���P��<P���    P��H                                                                                                                                                                                                        L       parents[$l#L       m���                                                           	   	   
   
                                                                                                                             !   !   "   "   #   #   $   $   %   %   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   :   :L       right_children[$l#L       m               
                                     "   $   &   (   *   ,   .   0   2��������   4   6   8   :   <   >   @   B   D   F   H����   J   L   N   P   R   T   V   X   Z����   \   ^   `   b   d   f   h   j����   l��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       m@��?�9X?�A.=q?�/@@  @kC�?�#?��D      D��    @�=qB�(�?��   >	7LB   B8  @ Q�@?;dD�`    Bg��F3=�D�3B���B�  B�\   @�ffA��@ Q�AP  B�     >@�Ǜp5      B�ffB�ff@��@@  D�  B4z�BY33�:$   @@  BR��         @fv�@�ffĝr�@�  �d��E��E��fŮ����[	E� 8��g�F�'I���rF��F�hS��(IƉ=�š�v�M�F�2�G8XNH��ZH��/{@E�AF��Ex��t�F�$�Cc6g��8��UK�KE�G �nE�tDr�4�v��Ƈ���ehg�8��.��EQ����A�ͻz�w&5F'�F��E����]��[�O�`y�F7W$ǅ<�Ŵ�L       split_indices[$l#L       m   	                  
                                             
   
                                        
                                                                                                                                                                                                                                                                                      L       
split_type[$U#L       m                                                                                                L       sum_hessian[$d#L       mF�` F�� CK  F� Cc  A�  C6  F�� C�  B�  B�  A�  @@  B�  B�  Fh� D�@ B�  Cj  A  B�  Bt  B\  @@  Ap  @   ?�  Bl  B   B�  @�  FV D�� D�` C�� B  B   Ch  @   @@  @�  B  B�  BH  A0  B4  A   @   ?�  A   @�  BD  A   A�  AP  Bh  A�  ?�  @@  FB� D�� D~� C$  Dz� C�� C�  @�  A�  A   A�  A   BD  C7  ?�  @   @   @�  B  @@  B8  A�  B,  @�  A   @@  B  A  @�  @@  ?�  ?�  ?�  @�  @   @�  Ap  B  @�  @�  A�  @�  @�  @�  B(  A�  @@  A�  @   ?�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       109L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       yA��E��*�+JF'��.1ň�~D(��GcE��Ŭ��Fpa3F\I���)ı�)E�gR�i�G+��ǝ��E�����R�GΩaG"�V��}�hN�F��/��t�FA�
D��
�ۀ�E����c��A�bƔ:�G��VF���F�AG���|E�\>Ǥb�GAp� ��G&��G��F�yOH VE���ZtEi���nP�H�F���ӊh�iyF߸��Ĕ�E.���W�D��i��}�jF�8`�Oy�ī��ƫ��k��E_KG �tFK��E���Gi�3�6��ōmmD��WF'����iǎT6E��!GnzD@�Ş#F���Ee�*��y�F*�|G�R�F�֬F����!��~E>ƢA�E��-��0~F#W5G��FF�#�ƓF�����L�7FS�ƂϬE�6�F��C��{���ù�E\x��Hm�ҫ�j^Nũ�oǟ����?�ħ9�E��v���	w,FXr�h��1!��y��L       
categories[$l#L       K                             	   
                                        	   
                      
                         	   
                                  	   
                                        	   
                         	   L       categories_nodes[$l#L                                ,   1   9   >L       categories_segments[$L#L                                                                *       8       E       FL       categories_sizes[$L#L                                                                                    L       default_left[$U#L       y                                                                                                         L       idiL       left_children[$l#L       y               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =����   ?   A   C����   E   G   I   K   M   O����   Q   S   U   W   Y   [   ]   _   a   c   e   g   i   k   m   o   q   s   u   w����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       yQJ�Q]NLQ�m�Q�F�Q��R�NQ�q	Q��Q��Q��Q�qKR$�\Q�4�QȢ8R,�QIN�Q�Qf��Qt\�Q��6Q�c+R ϨQL�QްNQ�kVQ�`�R9"Q��Q�zR�-�Q��    Px�Q�'�Q�?N    Q��Q�+4Qw6�QԺ�Q�~�O�L�    Q�o6Qԟ6QY��Q�BQ��R}�P��XQ��Q��bR��Q�(�Q�86Q�{mR$Q���Ro9�Rl��Q�H�Qk�Qڼ                                                                                                                                                                                                                                        L       parents[$l#L       y���                                                           	   	   
   
                                                                                                                                   !   !   "   "   $   $   %   %   &   &   '   '   (   (   )   )   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <   =   =   >   >L       right_children[$l#L       y               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >����   @   B   D����   F   H   J   L   N   P����   R   T   V   X   Z   \   ^   `   b   d   f   h   j   l   n   p   r   t   v   x����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       y         D�  ?��>uD�  D� <D��A33?2->o@�A  ?��T=�1   =��TB�  =t�   @�33B�(�>A�7@   ?]/@[C�   B�     B����A�b>�I�@   B�  F�AG>���B   BfffD�� BJ�D�� G��=�7L   @   @�  ?   ? �   =#�
>Xb?��?���>���>���D�    ?�yB.��@���D��    �k��E_KG �tFK��E���Gi�3�6��ōmmD��WF'����iǎT6E��!GnzD@�Ş#F���Ee�*��y�F*�|G�R�F�֬F����!��~E>ƢA�E��-��0~F#W5G��FF�#�ƓF�����L�7FS�ƂϬE�6�F��C��{���ù�E\x��Hm�ҫ�j^Nũ�oǟ����?�ħ9�E��v���	w,FXr�h��1!��y��L       split_indices[$l#L       y                                        
      
   	       	                        	   
                                                                        
       	               	                                                                                                                                                                                                                                                              L       
split_type[$U#L       y                                                                                                              L       sum_hessian[$d#L       yF�` E  Fg@ D�� D�  Ey  F(� C'  D�  DU� Cj  Cɀ E_� E҈ E~� A�  C  A  D�� DS� A   B�  C  C
  C�� EQ0 Cl  E�� E E< D�� @   A�  BX  B�  ?�  A   D�  @�  A�  DN@ @�  ?�  B�  A  C  Ap  B�  B  @�  C�  EJ0 B�  C%  B�  E� C�  E0 A�  D�` D�� D@  C�  A   A   A�  B   B�  @   @�  @@  D�� B�  @�  ?�  A�  @@  C�  C� @@  @�  @�  B�  @@  @�  A`  B�  A  @�  A`  B�  A�  A@  @   @�  A  Cy  D�  D�` A�  B�  C   B  AP  Bh  E D�  A�  C�� Dހ C� @�  A�  C�  D�  D�  C  A�  D9� CW  B�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       121L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       ]A�j�vF�%�D����F�>�G�}=ƄضD�/�F�B`�${*F������ŠRG�iD�V��,K�E�0�â�PG���wYŠ+3E
H*FH��GoV�E�d%��mF_��G�_F��ǫY-ƒ����~AF,O��a�F>8ĩN�H|�F������G��k���C�v�ŋ�tFzD��yGE�GɝF���Ft4�U�F��T'�t��7+nF�_�<�n�����?�QE�4Dn6�ăΙG#�E)z�F�� ĉ�TD���F�>G?�qDͭ�F�}wƭ2|�5��G�8Ä$�� ��j�El���P��
B��#4�E��A�2EFNd.�㯳F��|�'�@E;�G
*��+gF �Ŭ�gD�o�L       
categories[$l#L       *                                    	   
                                        	   
                                 
                L       categories_nodes[$l#L                         !   (   2L       categories_segments[$L#L                                                         (       )L       categories_sizes[$L#L                                                 
              L       default_left[$U#L       ]                                                                                L       idi L       left_children[$l#L       ]               	                        ����            !   #   %   '   )   +   -   /   1������������   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y����   [������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       ]QB`rQ:C�QE�Q�EDQ��Q�rPc�Q�q�Q��Q���Q���P� XP�t�    O�1PR&)AQ�1bQ��Q���R+ Q���Q�~�Q�~QP���P�#�O&��            Q�;Q�tQ���Q��R}�R�Q��8Q��OQ(HQv+�Q_�P?�LQ��R
ݢQ�b�R6�P��PS?�PPO"K�    N#�h                                                                                                                                                                        L       parents[$l#L       ]���                                                           	   	   
   
                                                                                                                 !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   2   2L       right_children[$l#L       ]               
                        ����             "   $   &   (   *   ,   .   0   2������������   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X   Z����   \������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       ]A�     ?   ?\)>���>;dZ@�     @B�\>�%?�M�>^5??ٙ�ŠRB8��>��^?!%?|�>C�   ?X��A�  >���>I�@�     ��mF_��G�_>���   @�  B�     ?���B�  @�  B z�C  @      A�  @@  A��>���<�B���B6ff>1'Ft4   F��T'�t��7+nF�_�<�n�����?�QE�4Dn6�ăΙG#�E)z�F�� ĉ�TD���F�>G?�qDͭ�F�}wƭ2|�5��G�8Ä$�� ��j�El���P��
B��#4�E��A�2EFNd.�㯳F��|�'�@E;�G
*��+gF �Ŭ�gD�o�L       split_indices[$l#L       ]                                    
                
             
                                                                                  	         	                                                                                                                                                                               L       
split_type[$U#L       ]                                                                                     L       sum_hessian[$d#L       ]F�` F�� Bd  Fd E�� B@  A  CX  F C  E�  B  A  ?�  A   C   B�  E7  E�x B�  BX  E�� E� A�  A`  @�  @@  @�  @�  B�  A�  Bx  A�  D�� Dk� D� E� A�  B�  BD  @�  E%  D�` D�  D�� A�  A   @�  A   @   @�  B�  A�  AP  @�  A�  B0  A@  A`  DS  D�  Dj  @�  C�� A�  E�@ D�  @�  A@  B�  A�  A�  A�  @�  ?�  E� C�  D%� D�� D�� B�  Cـ D$� @�  AP  @�  ?�  ?�  @�  @@  @�  @   @   L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       93L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       QA�:	B��Lƪ�.�:�E1֭Ǘ)��aV5É>ƒ-�F�ڽE�������^��2����F��kU;ƈBtń +�MN��8<�GW�E��.Ŋ5��M{�FC�k��a'�&$N��d�����HE1�]�GJ�F
����cmG�H�_F�,EL fCu��"nE��(@�F�|�^KB�X�F.��D��9�*2�D��=��F&��B<E5-���G�!qk4�݂��Z���F*�D����E�0�G	6�F��^G�2F�~F�_PE�#A�ݷG��;�A�x�Q��ħQ�D~���}f�D{FJa��z�ƪ�aL       
categories[$l#L                                           	                                L       categories_nodes[$l#L                         &   *   ,L       categories_segments[$L#L                                                                L       categories_sizes[$L#L                                                               L       default_left[$U#L       Q                                                                     L       idi!L       left_children[$l#L       Q               	                  ��������   ����               !   #   %   '   )   +   -   /   1   3   5   7   9����   ;   =   ?   A   C   E   G   I����   K   M   O������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       QP��Q\�P�=�Q�	<Q�)wOA=�P\��Q[�BRG�Q��Q���        PB`,    QF�JQ�TGR��Q��Q��[Q��R�Q��P�XP.�Q�mRh2�Q�_�Q�O�Q�aQ��Q�sx    Q�XP\��Q#t�Q��pR�QΟ�Q��Q�޼    O���O0��P��                                                                                                                                                L       parents[$l#L       Q���                                                           	   	   
   
                                                                                                               !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   *   *   +   +   ,   ,L       right_children[$l#L       Q               
                  ��������   ����                "   $   &   (   *   ,   .   0   2   4   6   8   :����   <   >   @   B   D   F   H   J����   L   N   P������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       Q@��;?"J>�\)?+C�=u   B�  ?5?Btp�>��?��������^�@   ��F�B�  B�  Bq33AP  @��      @�     @@  B�  ?��/   @   ?z��>��D�  GJ�=D��@@  ?9�B�  ?ȴ9   =#�
@�  E�   B<ff   B�X�F.��D��9�*2�D��=��F&��B<E5-���G�!qk4�݂��Z���F*�D����E�0�G	6�F��^G�2F�~F�_PE�#A�ݷG��;�A�x�Q��ħQ�D~���}f�D{FJa��z�ƪ�aL       split_indices[$l#L       Q   
                           	                                                                
                         
      	                                                                                                                                                                L       
split_type[$U#L       Q                                                                         L       sum_hessian[$d#L       QF�` F�� B�  FKd E�� @�  Bx  FF0 C�� B�  Ez� @   @�  Bt  ?�  FC  CD  Cj  B�  B  B�  E'� D�� A�  B0  F8| D*@ C7  AP  Ce  @�  B�  ?�  A�  @�  BT  A0  CO  E� D�@ Cr  @   Ap  A   B  F7� BX  C�  C[  B�  Bh  @�  A  B�  B�  @   @@  B<  BL  A@  A�  ?�  @�  B@  @�  A  @   C   B�  C�  D�  ?�  D�  B�  B�  @@  A@  @@  @�  B   @�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       81L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       UA�)�#�gDE֩�B�G?�bD;�Ga�w��7rƫ�G~����E�	�r�Q�BF�K�����ǧ��G��/�m���f���fG��2E(WG�_�R�  ��1�wE�ӁH�E5���)��nE���G@�zG�|ŖS�ưG�C�c��#0�"�G�2C����F^E�H �F��;EU��r7ä�g�	ЙD�>V��ME��t��?FG�MGz�(F]�S���>�Vm���/�ǭ)�F�k�Ť�%F��D�5�GD�sF%u��e8�^���������G*F&����@1E�F5�D�?�F�E�Gr��D���G{�D����h�rD����v'L       
categories[$l#L       6                                    	   
                                        	   
                	                           	   
                            
            L       categories_nodes[$l#L             
               !   "   &   '   (   *L       categories_segments[$L#L                                                                                             +L       categories_sizes[$L#L                                          	                                                 L       default_left[$U#L       U                                                                        L       idi"L       left_children[$l#L       U               	   ����                                 !   #����   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A������������   C   E   G   I   K   M   O   Q   S��������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       UQ�!Q���Q��Q�o�Q(�XQ�U�    Rl�Rq��Q.X�O�R�jQ��R+��R��R_edR�((P�GHN-?p    M��QI��Rb�Q�}�Q~��Q�),R9-yRX��R6��RGPQ�O�RX��P�`P�P��            J��N�c�Q�@Q��PRXj�Q�Q�60Qa7�Q�s�                                                                                                                                                        L       parents[$l#L       U���                                                     	   	   
   
                                                                                                                                   !   !   "   "   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .L       right_children[$l#L       U               
   ����                                  "   $����   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B������������   D   F   H   J   L   N   P   R   T��������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       U?��A@  C  B�     D�  Ga�wB�  >�A�     =u=<jB�  @�  @���B�  D�     �f�A�?��   =���   @��@@     @�H>2-A�  D�` >,1      ŖS�ưG�C�c�         D�     @�  A��?�p�?�M�ä�g�	ЙD�>V��ME��t��?FG�MGz�(F]�S���>�Vm���/�ǭ)�F�k�Ť�%F��D�5�GD�sF%u��e8�^���������G*F&����@1E�F5�D�?�F�E�Gr��D���G{�D����h�rD����v'L       split_indices[$l#L       U                                      
   	                                                                	                                              	                                                                                                                                                           L       
split_type[$U#L       U                                                                         L       sum_hessian[$d#L       UF�` Ep� FP� En� B  FP� @   E^� C�� A�  @�  EP� FL EQ� CP  CO  BH  A�  @   @   @�  A�  EO B�  F< EK@ B�  C4  A�  CB  AP  A�  A�  A�  A   ?�  ?�  ?�  @@  @@  A�  E� D}� A   Bp  E*� E�  ED� B�  B,  Bd  C!  A�  A@  A�  B�  B�  @�  A  A�  @�  @�  A`  Ap  @�  @�  @@  ?�  @   ?�  @   A�  A   D�� D{@ C�  D8@ @�  @@  BP  A   E� C]  E
  E�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       85L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       {A̵*�-x�EZ"f��O�s�.D�m�F����*3+F��N�#WDл �P�E��tGb��ƚ=�ݙƹ2hG�7�FzS�#�ǲ���
x8G�b��$�E^�REW6�Gc0�G�+rFt;�G0�^�MC{�M���C��G����jGFG�ZzG@*4�ÇD��dw��ځG0g�FM�/�P�G[�GF�[��qr���M�w]G�F��l��{�G�CHh/�G�CGO�H&E;��`��GĺǭIĜW9��Ô�1Z������5��s��G;��pXEF�F�/Z�oF	��G QgG=o(F :���~;D���<8EA:}āC���YqjƟD^�O�F����bЊƥ��F^�dƢH-ơ9F̢oF qq�"@xG%�"�_*F���<SE`�GGsΙB��?ƶ�|F��ŁdiF�I�G�%=Gag�F�ÃF�N��FNNgGMڋŠSoF��OF[ ���E���G+OR���]E��gFR ^�G��L       
categories[$l#L                                      
                                      	   
                     	L       categories_nodes[$l#L                   ,   8   ;L       categories_segments[$L#L                                                  L       categories_sizes[$L#L                                                 L       default_left[$U#L       {                                                                                                         L       idi#L       left_children[$l#L       {               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S����   U   W����   Y   [   ]   _   a   c   e   g   i   k   m   o   q   s   u   w   y������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       {Q�[Q/]�R�QnbTQ�X&Q� Rb��Q��cQۢQ��<Q���R359R�FQ��Q��"Q!eQ��GP��Q���P�(^R'�<Q�W�Q�"cR#�Q�D�Q�(�RH1�Qһ�Q�Q鿖Q��/Q��MQK�TQ��:Q�iyP���Ob1@Q�$�QO�P?WVP�Z�Q�\�    Q�'[Q�H    P�$Q�� Q�+�QdKQ�KR�+TQ��QsU�Pg Q�lHQ�R�N�ـQC Qu�xQ@�QApQ��                                                                                                                                                                                                                                                L       parents[$l#L       {���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   +   +   ,   ,   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <   =   =   >   >L       right_children[$l#L       {               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T����   V   X����   Z   \   ^   `   b   d   f   h   j   l   n   p   r   t   v   x   z������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       {?z�?��B�  ?�?b      ?�   Bg��B���?j=qA�  @"^5@���@@  =�Q�D�@ >W
=D�� ?o>��?�;>���A�H?L1E}  ?
��=u?�dZ?�bN><j?�n�A  @`B?H��A�
=?rn�>�%=�O�>��j>��-G0g�A@     G[�G@���?�7L?��=\)@�C�?G�B�  ?=p�B4z�@�     @��R@U�T   @XQ�@��?��!��Ô�1Z������5��s��G;��pXEF�F�/Z�oF	��G QgG=o(F :���~;D���<8EA:}āC���YqjƟD^�O�F����bЊƥ��F^�dƢH-ơ9F̢oF qq�"@xG%�"�_*F���<SE`�GGsΙB��?ƶ�|F��ŁdiF�I�G�%=Gag�F�ÃF�N��FNNgGMڋŠSoF��OF[ ���E���G+OR���]E��gFR ^�G��L       split_indices[$l#L       {   	   	      	   
         	             
                                 	         
               	               
                                         
         
      	                
             	                                                                                                                                                                                                                                                L       
split_type[$U#L       {                                                                                                                     L       sum_hessian[$d#L       {F�` F^� E8� F[L CP  E-� C3  FY< C  B�  B�  D&� E� B�  Bp  FW C  A�  B�  BH  B   B�  Ap  Ce  C�  E p B`  B�  B<  A�  B   C�  FR� A  C  A   A   A�  B�  B(  A   A�  @   B|  B@  @�  A0  B�  C   C�  B@  C�  D�` BL  @�  B   B   @@  B0  @�  AP  A�  A�  A  C}  FR( BH  @�  @�  B�  B0  @�  @�  ?�  A  @�  A�  @�  B�  A   B  @�  @�  A   A�  B<  A�  A�  A�  A  @   B�  @�  BX  B�  @   C�  B  A   C�  A   DĠ A`  B  A�  ?�  @�  AP  A�  Ap  A�  ?�  @   B  A0  @@  @�  @�  A   A�  @@  A   A  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       123L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       gB1�yD�6���>�E�;ŏ�U�E7�1~�Eg����ŧ8sHKy�E�F<C�Lk	H
��E��q�8�}Fp�Ž<����GN�#G��?F[��L��D2�F�̐���������nH5E��Et1�FE��Ƣ�CĄ�Gz΂F��ߵ�� w)F2^��"��Ǭ�G�~�Ā2G�-�밝ǂ'E@��GeňF�����ͪ��4� G**^�Z�FȞ�Gs>D�W$ŋ2�E��D�:�Ń���t��<�iE�C�GkE�DͯJF�˄D�-���ƁS6ņ��C�EX1GU]5E�Z�ň,��,3���G,��FC%�C�)�7ZG+�
�vĭ�
Ɔ���zD��"E��Ɯ+ G(�F��E\&iG4�F+�P�^� Ż��Ƽ����Ǉ�BMLl�6_�L       
categories[$l#L       +                             
                         	   
                                   	                                             L       categories_nodes[$l#L                       
                  -   3   4L       categories_segments[$L#L                                    
                                   !       "       #       %       *L       categories_sizes[$L#L                                                               	                                   L       default_left[$U#L       g                                                                                    L       idi$L       left_children[$l#L       g               	                                    !   #   %   '   )��������   +   -   /   1   3   5   7����   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c����   e������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       gQkVQRV�QlD;Q^=MRS�Q���R��R��Q��LQ��0P4�0Q�w�RPQ�PZ��Q��Q�WQǩQ�j�Q���R!��        Q�IhR/�RTX�Q�wQR4�vQu?�OF@@    Q���R�FQ�z�Q��R��aQ��R�`Q�"�R
q�Q���N���Qc XQ�&XQB.�Q���RJ��RTFR���Rk��Qu#Q��jQ010    Q>�T                                                                                                                                                                                                L       parents[$l#L       g���                                                           	   	   
   
                                                                                                                       !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   6   6L       right_children[$l#L       g               
                                     "   $   &   (   *��������   ,   .   0   2   4   6   8����   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d����   f������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       g   A�     @�
=>�1@陚B�        ?2-   @�        @ə�D�  >�$�?�^5?Z^5   D� G��?F[�@jn�D�� @   D�` B��D��    E��   >�K�B��{A�  @�  @أ�BZ  ><j>Ǯ>7K�B�RD�  @��D��    B�  B�  ?Z��B��{@�ff      G**^@�ffFȞ�Gs>D�W$ŋ2�E��D�:�Ń���t��<�iE�C�GkE�DͯJF�˄D�-���ƁS6ņ��C�EX1GU]5E�Z�ň,��,3���G,��FC%�C�)�7ZG+�
�vĭ�
Ɔ���zD��"E��Ɯ+ G(�F��E\&iG4�F+�P�^� Ż��Ƽ����Ǉ�BMLl�6_�L       split_indices[$l#L       g                                                     
                                                    
                                                 
                                                                                                                                                                                                                    L       
split_type[$U#L       g                                                                                          L       sum_hessian[$d#L       gF�` F� E�  F� D�� Eʘ D@ E� E  D�@ @�  E�� D]� D� @�  E� E  C�� D٠ D�� A�  @@  ?�  E�( D-� C�  D@ C\  Cŀ @�  ?�  E$� D�@ C\  E@ B  C�  Ch  D�� Co  D�� @�  A�  E�� A0  D@ Bh  C2  B�  C	  C�  CU  @�  @   CĀ @@  @   E` C�  D@ D�  CN  A`  D�� B�  A0  A�  A   C�  B�  B�  C D�  Ck  @�  C  Dx� @   @�  A   AP  Ew� Dh� @�  @�  D� B  B  A�  C  A�  B   B�  B�  AP  A�  Cр C@  A�  @   @�  C�� B  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       103L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       gBA 8�B�6CT��`drF�{��^	D(����H��G6�=�/8��`��¬F��fD�E�0�t�PrF:�.�E%�E���F�ZE������1�e�Fم���rdEi�F}�G���ã2�EW��Ƒ���sޜF�l��ؽLG	�E��d�vd�F���EAgÁ� E�A����hE���H.���B��Y�GCE5�LW�5Z�F��hG5��F�tD��ų�E��G"<@��͐Ec4Ƣz��?w4ě0Fc�Ű�r�x.�EWהFG<Ea�q�Z�AFatZţ�	FE���TJF ��]�C ��ìAE��f�@ԩGv��E��3ǌl���c�F�z��4WG,�F�DFP��Ɠ,��ָ���~F4���Ƽ�F���W-�D7�(Ĉ5D*$�š�JDp�_�:��F�Z���L       
categories[$l#L                                                                                                   L       categories_nodes[$l#L                
         *   4   6L       categories_segments[$L#L                                    	                            L       categories_sizes[$L#L                                                               L       default_left[$U#L       g                                                                               L       idi%L       left_children[$l#L       g               	                                    !   #   %��������   '����   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G��������   I   K   M   O   Q   S   U   W   Y   [����   ]   _   a   c   e����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       gQ��P��PܠdP� O�g�Q���Q-�P���PT��NG�NQb~Q��RL;dQ��bQ-�PH�|P�y�O���P=        LTp�    Q�u�R�,�Q��hQ�e�Q_�iQO��Q^��R��N�lO�z�P�-O��N)�@O55�P7�O�z(        Q�q�Q���Q�*xQ5(�Qu� Q���Q&�Qt6�P\��Q��"    P���Q��LR]�Q��~Q�>                                                                                                                                                                                        L       parents[$l#L       g���                                                           	   	   
   
                                                                                                                       !   !   "   "   #   #   $   $   %   %   &   &   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   4   4   5   5   6   6   7   7   8   8L       right_children[$l#L       g               
                                     "   $   &��������   (����   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H��������   J   L   N   P   R   T   V   X   Z   \����   ^   `   b   d   f����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       gA�  @U/=���   E}  D�� =�{>�   D��    ?>@�>�1D�     >}�>��wAp  E���F�Z   ���1>���B�  =ě�@R�\D� D�@ D�� A  >ȴ9A   @�  @   @�  ?���>�Q�BT  EAgÁ� >\   By33@�  @�  B�=q<�B(��>�{>��;G5��   @�     A�  >��/��͐Ec4Ƣz��?w4ě0Fc�Ű�r�x.�EWהFG<Ea�q�Z�AFatZţ�	FE���TJF ��]�C ��ìAE��f�@ԩGv��E��3ǌl���c�F�z��4WG,�F�DFP��Ɠ,��ָ���~F4���Ƽ�F���W-�D7�(Ĉ5D*$�š�JDp�_�:��F�Z���L       split_indices[$l#L       g                                      	                   
                      
                        	                                                         
                                                                                                                                                                                                                L       
split_type[$U#L       g                                                                                               L       sum_hessian[$d#L       gF�` C^  F�� CU  A  D�` Fl< B�  C  @�  @@  Dހ B�  B�  Fj� A�  B   A�  B�  @   @�  @   ?�  D�� B�  A�  BD  B�  A`  F4� EY@ AP  A�  A@  A�  @�  A�  B�  A  ?�  ?�  D@ D�� B�  A   A  A�  A�  A�  A`  BP  @�  A   F� D�` ER� B�  A@  ?�  A�  @   @�  @�  A�  @�  @   @�  A�  @�  @   B�  @�  @�  C  CĀ D+� C�  Bp  A�  A   @   @�  @   A   AP  @@  A�  @�  A�  @�  A   B<  @�  @@  @�  E� E7� D�` D2  EN B�  B�  B  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       103L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       sB�cį�(D�Ǖ�\.�����E�]�B2]9E��Ŋ�EP���4&�E�-���w�{Y�D��@F��|Dg�����*F�rŦ�qF��M�R���O�FOK�S����ǟ������P��Ɔ��D��F�HGD�V;��yŢ@�h��q�G�E�4Y��S�Ƹ6`Ƿ�HF���V'�*�F��[G37���s<�^g��_F�kƃQ�������E�2|�,Š�&EE���9��E��EF�,�G�>�C�»G�n� D�؊D�Ӟ�{��;"�n FC��z xG*`ĀO�F0��ąL�E��,�$0�Fң���o~�E��"D��*F!��F�J�E7�2�f1D�!�FƤ`F�	��g�Ŕ��Ɯ�
ŅJRƣ�ŘT��ϏFQ�Ƃ��N��v��Ɓ��E���ǖ�Ʀ��F�7h�2��Ɵ�`C�Wv���FgB��BE�L       
categories[$l#L       3                                      	   
                             
                      	   
            	                                           	   
      L       categories_nodes[$l#L                         %   (   /   0   2   7L       categories_segments[$L#L                                                                       !       #       'L       categories_sizes[$L#L                            	                                                        L       default_left[$U#L       s                                                                                             L       idi&L       left_children[$l#L       s               	                                    !   #   %   '��������   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c   e   g   i   k   m   o   q��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       sP�XQ�l:QK�$Q�YQ�)0Q�tXQ�?�R�:Q��|Q�OQ�erQ��Q?��R'ĞQ_�R@r6R��R8��RҩP7 �        Q�"lQ��Q\�sP�N�O�C@QӻQ�N�Q�2Qf`�R[�Q�_PR|~�R��DQ��R �nRxR�MrP�"PUQ��RKj[R	�rQ��KQJ2Q��4P6+O�њO��O�0 Q�-wQ�ǳQ���Q�ɠQ��>Q���Q͕�Qyy�                                                                                                                                                                                                                                L       parents[$l#L       s���                                                           	   	   
   
                                                                                                                             !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   :   :L       right_children[$l#L       s               
                                     "   $   &   (��������   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d   f   h   j   l   n   p   r��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       s?%�?"M�>�      D�  >2-D�  @�  ?a��D�     ?�ff>��m=��
?9XB�  D�� B���   F��M�R��B�  ?�l�@�     BI��>��B���?a%?3��=ȴ9B��=B�  B�  >F��>(��   B�  B2�\   =t�B��{?L1B�B�?'�@)�#      A     D�� Brff@�  >+   ?���A`  A   �9��E��EF�,�G�>�C�»G�n� D�؊D�Ӟ�{��;"�n FC��z xG*`ĀO�F0��ąL�E��,�$0�Fң���o~�E��"D��*F!��F�J�E7�2�f1D�!�FƤ`F�	��g�Ŕ��Ɯ�
ŅJRƣ�ŘT��ϏFQ�Ƃ��N��v��Ɓ��E���ǖ�Ʀ��F�7h�2��Ɵ�`C�Wv���FgB��BE�L       split_indices[$l#L       s   
   
                                            
                          
                                                              
                                           
                                                                                                                                                                                                                                      L       
split_type[$U#L       s                                                                                                        L       sum_hessian[$d#L       sF�` F x FH E�X C  D�� Eڨ E�� Ei� B@  B�  D�� B  C� E�p CC  E�p EL  C�  B4  @@  @�  B�  D~� Dg@ A�  A�  C�  B�  C*  E�  C/  A�  E{0 B�  EG� B�  C�  B�  A�  A�  B�  A�  D"  C�  DP� B�  @�  A�  A0  @�  B�  C�� B�  A�  B�  B�  D�� E�x @�  C+  A�  @@  EzP A`  A�  B�  D:@ E0 A�  BL  B�  C�� B  B�  @�  A�  @@  Ap  @   B�  A   A  C�� C�� C�� A�  Ct  D� B�  A�  @@  @   Ap  @   @@  A   ?�  @�  B�  AP  C`  B\  B|  A�  @�  AP  Ap  B`  BL  B@  D�@ B  ED� E  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       115L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       uA�� ����DX��8���`՝�D�bnEm��ŅۑƼ�F����ǨEpŪ�D��EYxKG܋UE+���,��E��E_W�H:A*��*+G-b.Fo)����`F�E��tE>����bF.��ß�NGn�GS��Ķ�QFl���e ��Ӥ��$�+G���ŹcOG���G4
�"�:HrӆFFy E6��e�tF�m��HZ��B����E��G�Pi�e�Ű}E��\ŠB��7�Ԭ�E �<F���FT�����oF�f�D �F:�u�@��4IF=�%��V�*[��R�CFG"��	O����ŬƧGF�/Ɯ�E���F�'���1����F�������sηG�����f4��;�F�!���F��E�B�Ʈ8�Cr �����E���E��a�+�����+�!E������Gf�h�1�5�T���F�H�D�/��\ ��r���j^TĎ��E����z�[ſ6�L       
categories[$l#L       ?                                        	   
                                         	   
                        
                                  	   
                               	               L       categories_nodes[$l#L       
                         "   #   3L       categories_segments[$L#L       
                                                          %       2       >L       categories_sizes[$L#L       
                            
                                          L       default_left[$U#L       u                                                                                                   L       idi'L       left_children[$l#L       u               	                                    !   #   %   '   )   +   -   /   1����   3   5   7   9   ;   =   ?����   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]����   _   a   c   e   g   i   k   m   o   q   s��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       uP�*�Q���Q��oQ�r�R>_QxyJQ9��Q�n�Q�4~R WR���Q�QOLNQ��Q\�kQ]�P���Qx��Rz��RYDQ�`Q�|�Q���P�#ZP��    Q#��R+��Q�X0Q�WQ�CQ�
�Q��0    O9Z�Q#�R/4&RncrR{=�RF��P���Ra1QY|�Q���Q��:Q��P&P#B�P��*    NF�O�P��(Q���R3A�Q�pQ��Qȶ�Q�O3R0�RI*�                                                                                                                                                                                                                                L       parents[$l#L       u���                                                           	   	   
   
                                                                                                                                   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <L       right_children[$l#L       u               
                                     "   $   &   (   *   ,   .   0   2����   4   6   8   :   <   >   @����   B   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^����   `   b   d   f   h   j   l   n   p   r   t��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       u      D�� D�  @�p�   @@  A�  @@  @�  @IG�@33A     A        BI��D�� C  B���D�` @�@@  >��Fo)�@@  A�  ?�(�   B�  @�  >�Q�Gn�      D�� B�  B�  B�  @�  ?)��>333B`\)B�(�@�  Ba��>��>7K�F�m�B<ff   =�G�>���B^��D�` B   A   B�  D�� D�� E �<F���FT�����oF�f�D �F:�u�@��4IF=�%��V�*[��R�CFG"��	O����ŬƧGF�/Ɯ�E���F�'���1����F�������sηG�����f4��;�F�!���F��E�B�Ʈ8�Cr �����E���E��a�+�����+�!E������Gf�h�1�5�T���F�H�D�/��\ ��r���j^TĎ��E����z�[ſ6�L       split_indices[$l#L       u                                                                                                                                                                                                                                                                                                                                                                                                                                  L       
split_type[$U#L       u                                                                                                           L       sum_hessian[$d#L       uF�` E�� F<� E�@ C� BH  F< D�� E#0 C�� B�  B  A�  D�` F+@ D�  @�  D�� D�� C�  B�  B�  A0  A�  A  @   Ap  C+  Db  E�� E3� D'� D�@ ?�  @�  Dn� C�� B�  D�@ C|  @�  B�  A�  B(  A�  A   @@  A0  AP  @�  @�  @�  A0  C  A�  B�  DE� E�� Dw  E(� C,  D@ B  B  D�� @@  ?�  A�  Dh� C*  C  B�  A�  D�� B�  CT  B   ?�  @@  A�  B�  Ap  @�  A�  A�  A�  @   @�  ?�  @   ?�  @�  @�  @   A0  @   @   @   @   @�  @�  A�  B�  A   A   B�  A   D@@ A�  Eܘ B   Dm@ B  E� C�  @�  C'  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       117L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       uA<��ŝawC�΍��S�E�qÔ��EgU�D\���,V�C؂�G!�sAO�Ʋ��D���Fkk^���F+M�ſ�(ƈ8|�s�G<��EK#�GցDkņD����j� GmFD1�^EN�Gsu`DYL��i��F��`�U�oQ�EvJK���D��0SE%mƾsVG���^��E�u���  Ĭ�hE8`�FH��j��j�G���F�#�ǲ��Hh��MG���C�*�Ł�vG`��H�?F�������E�Lƞ���d���p\E��nDi���U ���o������FFnÔo���E%W�ٟ�C�Z�FY��E�)X�'@zF�QDE�&�C��ŕ�4�//�E��C�RE��D��pF��B���ť�ZD�
��-EG*+��I���
�WF�N�$�E�կGw!�E&���>*�F�MG>���M6�Ř�HD]�D��?�L�7G'�o��F���Gr"��ш^FKs�L       
categories[$l#L       7                           
                                             
                                                                  	   
                         	   
   L       categories_nodes[$l#L                               #   (   ,   2   5   7   9L       categories_segments[$L#L                             	                                                 !       #       $       0       1L       categories_sizes[$L#L                                                                                                         L       default_left[$U#L       u                                                                                            L       idi(L       left_children[$l#L       u               	                                    !   #   %   '   )   +����   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q��������   S   U   W   Y   [   ]   _   a   c   e   g   i   k   m   o   q   s��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       uP��P��`Q �IP��P��;Q��Q��P��[P�n�Pu�)P�rQG�dQ���Q��ARi��P��P�|�Pِ~P��8P��MP3<N��    Q?��RA� Q�Q�*vR�QH��R	RS��PKu�P Y|PHP8��P�I�P�$Pu� P�j�Pm��PV9�N#׀        M�AQ��vQ�e�Q>m�R�tQa�JQ	�pQe��Qɭ�Q�(Oӏ�P���QOo�QɻyRv��Q�k|Q��                                                                                                                                                                                                                                L       parents[$l#L       u���                                                           	   	   
   
                                                                                                                                   !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <L       right_children[$l#L       u               
                                     "   $   &   (   *   ,����   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R��������   T   V   X   Z   \   ^   `   b   d   f   h   j   l   n   p   r   t��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       u@   A   ?�   B�
?o@�  @3�
@�D�� A�     B���=u>�5?   ?�/>���>�JD�     D�� GցA�  B\)Bz=q   @@  =�w?z�      ?   =oD��    B   ? ĜA�  D��    A�  �^��E�u�   B���>�9X>�+?j=qB@��   D�  D��    Brff   >gl�   ?���D�  ?�!����E�Lƞ���d���p\E��nDi���U ���o������FFnÔo���E%W�ٟ�C�Z�FY��E�)X�'@zF�QDE�&�C��ŕ�4�//�E��C�RE��D��pF��B���ť�ZD�
��-EG*+��I���
�WF�N�$�E�կGw!�E&���>*�F�MG>���M6�Ř�HD]�D��?�L�7G'�o��F���Gr"��ш^FKs�L       split_indices[$l#L       u                                                                                               	                                                                                               
      
                                                                                                                                                                                                                                L       
split_type[$U#L       u                                                                                                       L       sum_hessian[$d#L       uF�` D�  F|` DF� C~  FT4 E � Cr  D
  Cs  A0  FQX C7  E� C� C  B�  C�  Cn  Cm  @�  A   @@  F,H E@ C  B@  A�  EP C�  B�  B�  B�  B�  A�  C$  C  C   B�  CN  A�  @�  @   @@  @�  E�� E�� C�  D�  C  @�  AP  B  A   A  @@  E  C�� B,  A�  B�  A�  Bp  @   Bx  @@  B�  Ap  @�  B�  B�  C  A�  A�  B�  Bh  BP  CG  @�  @�  A�  @@  ?�  @@  @   E�h C�� E�� C̀ Cf  C.  D{@ Dp� B�  B|  @�  @   A   @�  A�  A�  @�  @�  A   ?�  @   ?�  C4  D�� C�� B`  A�  A�  A   A@  @�  Bx  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       117L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       3A�D�@ۡGn�B-�t�7���"��G�h�C���ܾX�]RƊ�KƏ��ø`�G$�=FKm�A�F|F����K�Ŧq��aj�Ɓi�(����3Gū�/C��<F�f��J��'�ƃ����xG�Nƹ��F��w���F�gB��ƶ�1G �E�c����ǀ\�ƨw:�{��F���M�E�Ŗ�F����ϚE��m�HL       
categories[$l#L                                 L       categories_nodes[$l#L          	                  L       categories_segments[$L#L                                                         L       categories_sizes[$L#L                                                        L       default_left[$U#L       3                                            L       idi)L       left_children[$l#L       3               	                  ����������������            ��������   ����   !   #   %   '   )   +   -   /����   1������������������������������������������������������������������������L       loss_changes[$d#L       3P��PQzQ#�PƜ�Q��O	Omc�QmJ�Q�#zO�D�P��4                P޷%Q��
Q�@Q�O;        P�E4    Qv�bQ�R�Q.(O�� O� �Qwq�Q��    O���                                                                        L       parents[$l#L       3���                                                           	   	   
   
                                                                                      L       right_children[$l#L       3               
                  ����������������            ��������    ����   "   $   &   (   *   ,   .   0����   2������������������������������������������������������������������������L       split_conditions[$d#L       3CJ  CB  D�@ @�  =#�
B�33B�  B�  =49X   >_;dƏ��ø`�G$�=FKm�?=p�A`     A,���aj�ƁiD�@ ��3G?Η�C              ?��   ƹ��CG  ���F�gB��ƶ�1G �E�c����ǀ\�ƨw:�{��F���M�E�Ŗ�F����ϚE��m�HL       split_indices[$l#L       3               	                  	                                              
                                                                                                       L       
split_type[$U#L       3                                            L       sum_hessian[$d#L       3F�` F�T @�  F�4 A�  @   @�  F�6 C�� @@  AP  ?�  ?�  @   @   F�b Cj  @�  C�  ?�  @   A@  ?�  Dg  FrT Ce  @�  @�  @@  C�� AP  @   A   De� @�  Fr< @�  A  C\  @@  @   @   @   ?�  @   C0  C�� A   @@  A  ?�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       51L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       m@�IE9�j��tE�4G<���H`�D�F�`ß�UG���F}1�E�8�Ŧ�,ŬA�D�2Rĺ�F�&
ǰ�C�K�G�F_�:���F��xE�'�9s�D���Fx�����ĈcEkzF3b�Ǝ?���NF�ڏ��O��Ȼ�5.D���j��6��{.G;SF���M�hu�Ƿ���Y�F_�7ǣ�� D�E���G���ƇNC��]���K�Q�E_9uG���D+�pF�9�D�s@�T<Ə\�DP~BE� �F��.�y��_�Eu����O�+��D���Dԇg��]�D�}gFv݅E /<GT��C:F�4�F��ŗX8�����E���96��ć�;Fc�$E�4��E߲}�I�sF��维G[Q)F�}��c'cƱe+�<G���j��Eo����Ca�D���ϛ�GC_ƅ�L       
categories[$l#L       #                                      	   
                            
                                         L       categories_nodes[$l#L       	                   %   )   8   :L       categories_segments[$L#L       	                                                         !       "L       categories_sizes[$L#L       	                            
                                   L       default_left[$U#L       m                                                                                                  L       idi*L       left_children[$l#L       m               	                                    !   #   %��������   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A����   C   E   G��������   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c   e   g   i   k��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       mP���Q)�bQG�Q)Q�Q

Q+��Q�|�Q�y�Q9RP%i�Q�H�Q�H�QE�`QTN�Q��pQ�C2O� Qz%�        N3r�P
�QY�sQ[�Q��R,X�Q��3Q�'Q�Q���R�Q݉nQ;^Q�.    Oj��Q�@Q?�V        N_��N��Ra;nQ(݌P<ëP��Q��R��RR
�eQ u�P��PR7oQ��P�S�Q��Q���Q�ѥ                                                                                                                                                                                                        L       parents[$l#L       m���                                                           	   	   
   
                                                                                                                             !   !   "   "   $   $   %   %   &   &   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   :   :L       right_children[$l#L       m               
                                     "   $   &��������   (   *   ,   .   0   2   4   6   8   :   <   >   @   B����   D   F   H��������   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d   f   h   j   l��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       m   A�     >7K�      >���>t�<uD�� ?��RB�ff>���>�BP  D�� ?�>�  >A�7G�F_�:   @@  ?��>���B�  >ؓuB�B�?;d<�9XC  >�+@@  >@�B�=q��O�>�x�   >-V�j��6�   D�� ?��D@p��D� CW
B�ff>�JB9��=�l�>p��@�  B�  Bl  A      @Co   D+�pF�9�D�s@�T<Ə\�DP~BE� �F��.�y��_�Eu����O�+��D���Dԇg��]�D�}gFv݅E /<GT��C:F�4�F��ŗX8�����E���96��ć�;Fc�$E�4��E߲}�I�sF��维G[Q)F�}��c'cƱe+�<G���j��Eo����Ca�D���ϛ�GC_ƅ�L       split_indices[$l#L       m                                         
                                             
      
               	                                   	                        
                                                                                                                                                                                                                             L       
split_type[$U#L       m                                                                                                    L       sum_hessian[$d#L       mF�` E  Fg@ E� A�  Ey  F(� DC  D�� @�  A`  DO� EE@ D�` FL C�  C�  A   DƠ ?�  @�  @@  A0  DH� A�  D�� D� B�  D�` E�� E�� Cp  C:  B  C�  @   A   BT  D�  ?�  @   @@  A   D?  B  Ap  AP  DW  C� B   D� B�  @�  C� D� B  E�� E�h A  CS  A�  B�  B�  A�  A�  C�� B4  @�  @@  A�  A�  C�  D�� ?�  @   ?�  @�  D=@ @�  B  @@  @   AP  A   @@  DT@ A0  C�  C  A  A�  C  D�  A�  B�  @@  @�  C�  B  D	@ A  A�  A0  D�@ Eo� Eq� D=  @�  @@  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       109L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       {A'�kD�}�X�iE�učdF*�Eĸ��D�+F���aQD�DG�{E�T��Y�C{2��{E���G2�9E�G�!.lG��P�-E��Gډ ���K�eB
G�VƜ��8rD��������Wܟ�y�G�*E�'�Gq��ƎV�G�)hD+�X��	������H!�rE���?^VF�X�EGc�F� H�L�Q\F��.��N�1G�!F��b�e%Ş@GE����t9C�3�FXqs��PE5�7�D���(�DI��G�5F0i�G$�.F�C��TF����k���{�F��Fk�GQ޼ǐިD��8�E�0�r�<FS����'E�GuGnnCE�;4C��_F<#�]��L�;G`��E�P�E�jC#�F��ƞ��GM~��N �W��b�xF��� 2��0WJG=JF ���`չE����<����ؤF ����&qF6C�F�ZšOBbdE�ĠE�Ztŧ�ašH����hG��C�A
L       
categories[$l#L       +                         	   
                                                        	   
                                              L       categories_nodes[$l#L                                7L       categories_segments[$L#L                      
                                    !       $L       categories_sizes[$L#L              
                                                 L       default_left[$U#L       {                                                                                                               L       idi+L       left_children[$l#L       {               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a��������   c   e   g   i   k   m   o   q   s   u   w   y������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       {P�G�Q�C.Q���Q��Q�S�Q狎Q��Q���RR6fQ��Q�Z�Q�mtR��Q��QS�!Qܑ�Q�ҟRFhRjeQ���R@�&Q��"Q�o�Q�,�O�)RLÇQ�*|Qى�R4
6Qu	�RV�QjۤR]�"Qi��Q�LUR�/bR�DQ���Q�,QMqCQ���Q�AQ'�Q�Q�-pR4��Qj�tP��QPܝ         O���R-X�Qā4Q���Q���R.`zRj�Q�`tQ�R��RO��R�w                                                                                                                                                                                                                                                L       parents[$l#L       {���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   3   3   4   4   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <   =   =   >   >L       right_children[$l#L       {               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b��������   d   f   h   j   l   n   p   r   t   v   x   z������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       {@B�\@@  D�� B�=q>��>$�?yX>��   B�  @�  >\(�@�     B�ffB}��>���?U=L��B���         D�`    =o=�\)@�  >���B�  >j~�@ ��   >�Q�=��#?\�@�>y�#<�h>�`B?�y>A�7B�  B�  D�  >(��?�RB��B(  �Q\F�B`  @S�
=��@�Q�   >�=qD�  =uA�  ?D�>O�;=<j�D���(�DI��G�5F0i�G$�.F�C��TF����k���{�F��Fk�GQ޼ǐިD��8�E�0�r�<FS����'E�GuGnnCE�;4C��_F<#�]��L�;G`��E�P�E�jC#�F��ƞ��GM~��N �W��b�xF��� 2��0WJG=JF ���`չE����<����ؤF ����&qF6C�F�ZšOBbdE�ĠE�Ztŧ�ašH����hG��C�A
L       split_indices[$l#L       {                  
                                                                                              
                                                                        
            	                                                                                                                                                                                                                                                L       
split_type[$U#L       {                                                                                                                   L       sum_hessian[$d#L       {F�` E�P F* E  E~� D� F!� D�  D @ Dv� E@� A�  C�� E� E�� D2@ D^  CL  Cڀ Dn@ B  D�� D�� A�  @�  C�� C  D  D�@ EҘ D�� D*  B  A�  DV� C#  B$  A�  C�  DT@ B�  A�  A   DW@ DB@ CC  D�� @�  A@  @�  ?�  @�  C�� A`  C  C�� C�� D�� D.� E�x C�  C�� D?  D)  @�  A�  A@  A�  A   B�  D7� B�  B  A�  A�  A�  A   ?�  C̀ D9  B�  B�  AP  @�  A�  @�  @   DD� B�  D&� B�  @�  C=  C  D�� @�  @   A0  ?�  ?�  @�  B$  C�  @@  A0  B�  Ap  A�  Co  C  B�  D�` C4  @�  D-� E¨ B�  C�� B�  C�� BP  A   D=  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       123L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       SA|^��O�F�d�D(&��YG�>�F(�BjܰFM�T�@ƺ	uE�0ZG\� �F�"��TC6�LG�D���ĜXG�߹��FŇ��h"gC��G8�"��Ǉ�qE:fZ�D�9F���H�KFD]�I�XD/�=�R��HE��F�8 F��}�>��G�?��� E�g�1�FX�E��pDU`z�.z�� ���%��D��A��U��ҩC3��Ņ��Fa�F�d{G��EP��G��]D��Q� ����C� J�L�s�gG�6�F'WFs�����`F�B'ŘS��P���F; G+�EY�����aĆ>ZA�@ ÷gE��L       
categories[$l#L                                              L       categories_nodes[$l#L                      %   'L       categories_segments[$L#L                                           	       
L       categories_sizes[$L#L                                                 L       default_left[$U#L       S                                                                          L       idi,L       left_children[$l#L       S               	                  ��������                  !   #   %   '   )��������   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M����   O����   Q������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       SP���P��P���QChyQ�?�Of��P]yQO�R�aQ���Q�X        M��pO_��Q�kQbRRNF�Q��7Q���Q���Q�Q���        M�O��P }Q�lQ�&�Q�~�Q̖�Q��PQ��Q���Q��sQƔ�P��Q)V)P���Q�?@P�O�QD�
    K*	L    M��                                                                                                                                                L       parents[$l#L       S���                                                           	   	   
   
                                                                                                                 !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   ,   ,   .   .L       right_children[$l#L       S               
                  ��������                   "   $   &   (   *��������   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N����   P����   R������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       SA�  A�  AP  A�  ?���B8��   ?\)@   >��T>��/E�0ZG\      >�Z@B�\D��    Ap  >hr�=���>��Ň��h"gA�  A�  BY33?�9@�  ?|�BY33>n��?�u>�;d=49XC     >���   B��3D�  A0  E�gB���FX�B�33DU`z�.z�� ���%��D��A��U��ҩC3��Ņ��Fa�F�d{G��EP��G��]D��Q� ����C� J�L�s�gG�6�F'WFs�����`F�B'ŘS��P���F; G+�EY�����aĆ>ZA�@ ÷gE��L       split_indices[$l#L       S                                                                                                           
               	                                                                                                                                                                          L       
split_type[$U#L       S                                                                             L       sum_hessian[$d#L       SF�` F�8 A�  FZp EH  @�  A�  FN� D8� E:� CT  ?�  @@  @@  AP  B<  FN( C  D� E9� A�  C  Bh  @   ?�  @�  A   A�  A�  ET  F( B�  A�  C�� C|  E @ C�  @@  AP  A�  C  A0  B<  ?�  @�  @�  @@  A�  A  @�  AP  EN  B�  D�@ E�� B8  B�  A0  @�  C�  ?�  C  B�  B�  E� Cǀ A  @   ?�  A0  @   A0  A0  B�  B   @�  @�  B$  @�  @@  ?�  @   ?�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       83L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       %A���@^��Gz[�B%rV�š�n��F�~	�J�F��V���P�/vA��KǉQ�GC�Q�!��HČ�H�Z���Ʊ���2�G�|Žd�ƶM�Ɓ%G��ƍ��F8����PmC���G�#Ř{g�t��F���G>O�E���*�F�DL       
categories[$l#L          L       categories_nodes[$l#L          	L       categories_segments[$L#L               L       categories_sizes[$L#L              L       default_left[$U#L       %                                     L       idi-L       left_children[$l#L       %               	��������                     ������������   ����      ��������      !����   #����������������������������������������L       loss_changes[$d#L       %P���P�<&P��@P��,Q�        P�/�Q�j4P(0P� P��M�ƀQ�i�            P>`    P��IP��A        Q6�Q���    O.�                                        L       parents[$l#L       %���                                               	   	   
   
                                                      L       right_children[$l#L       %               
��������                     ������������   ����      ��������       "����   $����������������������������������������L       split_conditions[$d#L       %CP  CB  D�` C&  =#�
�n��F�~	C  @�     >�C  D�` D�` �!��HČ�H�ZD�@ Ʊ��?��B�\Žd�ƶM�B�  B�  ƍ��?���PmC���G�#Ř{g�t��F���G>O�E���*�F�DL       split_indices[$l#L       %               	                    	                               
                        
                                        L       
split_type[$U#L       %                                    L       sum_hessian[$d#L       %F�` F�X @�  F�4 A�  ?�  @@  F�� A�  @@  Ap  F�� @�  A�  @@  ?�  @   A`  ?�  F�� @@  ?�  @@  A   Ap  @   A@  E� F%P @   ?�  A   @   @�  A   A   @�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       37L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       {AJ�ZC��+�?ET�w��E��F�e���aAV�:��ԻC�S$G	��Gaeœ|�����*P%D��xj���!���+<G�R�Ŀz��1�Gg\F��H1>ƃ|!GE.�Ƽ;Y� t�G�1ŜaCAF��g�	d���3��XXF�M��9ތ�B��G��ƔŰ����E4��GG���C�G��œ@ń��GI<�HLK�Gx�	E�Zf�z��G��W��F��Nj���yǈd�ǳ��Gun�Z��F����BPEݾ���E�AGy���q��H�D����Q(ƃ�-�X�=Fp����*ƍ�Ăz�G26Fr'��4��B�ng�2����G)�De�Gf'�E°�Db9��S|GƴE��@G�\���ES"��G�G� E���G��NE�H���5^GF��ĉ�C�0w�ǔ{]E�{%F�#8E�PM����F:|ơJ�G�yŀ���P�z�EVF>��G=���m��k�DZmGUj�ũ8 D2ML       
categories[$l#L       <                     	   
                         	   
                                  	   
                                                                 	   
                            L       categories_nodes[$l#L       	               "   '   )   :   ;L       categories_segments[$L#L       	               
                     !       (       5       9       ;L       categories_sizes[$L#L       	       
                                                        L       default_left[$U#L       {                                                                                                          L       idi.L       left_children[$l#L       {               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I����   K   M   O   Q   S   U   W   Y   [   ]   _   a   c   e   g   i   k   m   o����   q   s   u   w   y������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       {P�r�Q.h!R��P��R"��RK!�R��P�?Q�U�Q͵7R<%R�Y?Q��R>m�Q�~uRJ�Q�LbP��EP�}�Q���Q���Q��R��Q;V�R6�Q��$P��Q�UJP��RsrQ�^�Q=τQ�.�Q��Q��O�{ P�^    O|0P~� OQڣQ���Q���QɻR'��Q�rP�rBQ�OPʾ�R@Q?ddR�,Px�O�t�Q�A�R#F�    O, 0Q�P��R��Q�B�                                                                                                                                                                                                                                                L       parents[$l#L       {���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   $   $   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   :   :   ;   ;   <   <   =   =   >   >L       right_children[$l#L       {               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J����   L   N   P   R   T   V   X   Z   \   ^   `   b   d   f   h   j   l   n   p����   r   t   v   x   z������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       {D�� D�` >7K�AR{B�\)   >��@.v�Btp�=�E�?�bNB�G�A   B��>���@'�@3o@�  >y�#?���?�>��`   B0  >߾wB���   >�>e`BA  >�   B���B�     >�1A0  �9ތB�     >)��   >��>�%?W�P@�=��@�  B<ffA   D�� =�j>�ȴA�  A�  >Y�>ȴ9ǈd�      >�oB��q?3�FEݾ���E�AGy���q��H�D����Q(ƃ�-�X�=Fp����*ƍ�Ăz�G26Fr'��4��B�ng�2����G)�De�Gf'�E°�Db9��S|GƴE��@G�\���ES"��G�G� E���G��NE�H���5^GF��ĉ�C�0w�ǔ{]E�{%F�#8E�PM����F:|ơJ�G�yŀ���P�z�EVF>��G=���m��k�DZmGUj�ũ8 D2ML       split_indices[$l#L       {         	                                                    
      
                    	   	                                                        
                              
   	                                                                                                                                                                                                                                                                    L       
split_type[$U#L       {                                                                                                                  L       sum_hessian[$d#L       {F�` Fp� D�� Fb� D`@ Cd  D�` Fb B  D3� C3  B�  C  CZ  D�  FE� D� A�  A   A�  D/� Bt  B�  B�  A�  B�  A�  CP  A   B�  D�` FCh C  B�  D�  A@  A�  @�  @�  A0  @�  B�  D  A�  B0  B�  A�  B   A�  Ap  A�  B�  B  A�  @�  B�  B�  @�  @�  B`  A`  B�  D�� DK� F6� C  @�  B�  A   D7@ Dq  @�  @�  A0  @�  @@  ?�  @�  @�  @   @@  B�  A�  @�  D  @   Ap  A�  A�  Bp  A�  @�  A�  A�  A0  @�  A�  A`  ?�  @�  A@  @�  B�  A�  @@  @@  AP  @   @�  A`  B�  A  B�  @@  @@  B0  A@  @�  A   B�  A   D	� D@ L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       123L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       sA���Ă��DQ���M�1�zEKD����GA�6�~g��\GS�E�$Cv�PG�	�� ����G�d)E�[����D����u�G�D�EК%C���F�LEE%��3Q�G|�JF7j�E̋�Ɗ�`�Y��ƅ�iZUH
�*F����(q�|���w��F���D��D��hƓEF4 �G�u�G�:��
i���D��_�!�G%9E�^��4�ņ�F-�E�K2�� B�OMG(|���O�1�ED�[gŬ>�E��N��֚Fs:�GK��Fl��DE)���`D�����_�K���E�EFZ��
�,A���E��D��*�\r���H��j��F�ţ��3zF1�G�DL�F��N�n5�U�t���a�Q�*F ������8��E<�F���D ��C�w�Eb�M����CF���*fj��r
D�ܵF�N��S�E��8F�W�@�FU%F������^�В'L       
categories[$l#L       4                                         	   
                                  	                                                                           
         L       categories_nodes[$l#L                                            !   ,   /   2   <L       categories_segments[$L#L                                                                               !       "       %       '       (       *       3L       categories_sizes[$L#L                                   
              	                                                               	       L       default_left[$U#L       s                                                                                        L       idi/L       left_children[$l#L       s               	                                    !   #   %   '   )   +   -   /   1   3   5����   7   9   ;   =����   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c   e   g   i��������   k   m   o   q������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       sP`
Q��'QW�aQ�F1Q�Qu/�Q��Q��Q�Q��wQ*s�R¾QT��Q���Q�+=P��Q���Q�Q�<rQ��Q�SP�3�QW(Q�b$R��Q�A�Qv�    M�8�Qo1Qҭ3Ng]8    Oo��P��Q%URPk
UR�2Q��~Q�QI��P�tQ��"P -P�-�O��PiyBQ �Q��VQ��	R|i�Q��nQ�("Q�|Q��U        P�,1P���Q���Q��                                                                                                                                                                                                                        L       parents[$l#L       s���                                                           	   	   
   
                                                                                                                           !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   9   9   :   :   ;   ;   <   <L       right_children[$l#L       s               
                                     "   $   &   (   *   ,   .   0   2   4   6����   8   :   <   >����   @   B   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d   f   h   j��������   l   n   p   r������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       s   =49X   <oB�  D�  =#�
@@     D�� >�V>��            ?��@@  >	7L@      B#
=   <�@�  ?���?�(�G|�J   B�33Bv{   �ƅ   D�  >D��?ƨB�\)>��7?D�D�  ?9�@�  D�`    <�@      =�o@      @`B@��@Ϯ@kC�E�K2�� ?Ͼw@���D��    D�[gŬ>�E��N��֚Fs:�GK��Fl��DE)���`D�����_�K���E�EFZ��
�,A���E��D��*�\r���H��j��F�ţ��3zF1�G�DL�F��N�n5�U�t���a�Q�*F ������8��E<�F���D ��C�w�Eb�M����CF���*fj��r
D�ܵF�N��S�E��8F�W�@�FU%F������^�В'L       split_indices[$l#L       s                     	                                        	                	                                         	   
                           	                       
      
                                                                                                                                                                                                                                            L       
split_type[$U#L       s                                                                                                   L       sum_hessian[$d#L       sF�` E�H F� C� E�� F� D@ A�  C�  E�� B  D�� E�� @�  D� @�  A`  C#  C�� E�� D�  A�  AP  Dw� D� E�  EOP @   @�  C-  C�  @�  @   @�  A  B�  B�  B�  CL  B�  E� D3  D@ @�  A�  @�  A   @�  Dv@ CD  C�  Ei� D  E<@ C�� @@  ?�  C  A�  C�  B�  @   @@  @   @@  @@  @�  A�  B\  B$  B  B4  A�  C(  B  B|  A�  E�( C<  D  C  C�  C+  @   @@  @�  A@  ?�  @�  ?�  @�  @@  @@  B�  D]� B0  C  C=  C  E$� D�  Ci  C�� E'� C�  C�  A�  B�  Bd  A�  @�  C�  A   B   B�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       115L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       {A�TD9��Ğ��DЛ��l�ŷ�SE��D
oEڟGE<Ƴ����Eu�NGC�D�E���ǢEkq%F�DE��E� Q��6����E�LŔ�c��l�F�����Fs�G��\E��@���\Ŝ`%EtxF��1E�GB����Gk5�C��E=��G�L�F�Ժ�ߣ�^���,/OE����݉ů�G�S	Ƃ�-�{�dFn4
�!�G'nU�0���hܚGhr:H9���W� B�DF&9�ı����X��Ŕ>U�P6�E^[�F�����6��i�D��zEV'F�r����x��D�EG�mņb�D��C@��F�B�G���E�K�@�E��"�B���;��F"���[SFL��DnE�C��LƉ�G>�0�BLD���ƹ{zE!$�F'2�D+G�Ʋl�F�Z��ΛeG !E �VƑ�E"�ƙ9ī��G�QEp�TG�#QFFQ'Ƹ%�E�V��y�ÄX�E��G�/��EMR��l��z� L       
categories[$l#L                    
                                        	   
                       L       categories_nodes[$l#L                      &   -   1   6L       categories_segments[$L#L                                                                L       categories_sizes[$L#L                                                               L       default_left[$U#L       {                                                                                                              L       idi0L       left_children[$l#L       {               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q����   S   U   W   Y����   [   ]   _   a   c   e   g   i   k   m   o   q   s   u   w   y������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       {Po��Q�Q�gQ_V�R�vQ��RQ��QQg�bRw0Q40�QZ��R��R�R
sQ��Qx�LQ�$�R��iR
ϣQ�4�P�p�Q��lQ%�gR��RsLR�nR+�QO�RP&Q�d�Q�Q��Q��R��Q�3�R2Q�E�RuQ�&�Q��R<��    P�b:Q�PQ�Pt�    Q}#^Q�jR.�dQ�j8R�=RC��Q�~Q�:P�(-Q���Q�mP�
*QdRQ���Qc��RP�B                                                                                                                                                                                                                                                L       parents[$l#L       {���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   *   *   +   +   ,   ,   -   -   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <   =   =   >   >L       right_children[$l#L       {               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R����   T   V   X   Z����   \   ^   `   b   d   f   h   j   l   n   p   r   t   v   x   z������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       {@��@I�?��y@��R   A��?��m?�!>��D�� ?���B�  D��       D�     >�+D�  D�  =#�
>��@�  B~=q?��B��>�>��?��RBl  B�  >��\>�l�@�  >+BD  ?���Brff   @���>�F�Ժ@@  ?T9X@      ��݉=�%@�     >>W
=@@  ?��   >k�A   B$  >��>��;>�?}D�@ ?j=q��Ŕ>U�P6�E^[�F�����6��i�D��zEV'F�r����x��D�EG�mņb�D��C@��F�B�G���E�K�@�E��"�B���;��F"���[SFL��DnE�C��LƉ�G>�0�BLD���ƹ{zE!$�F'2�D+G�Ʋl�F�Z��ΛeG !E �VƑ�E"�ƙ9ī��G�QEp�TG�#QFFQ'Ƹ%�E�V��y�ÄX�E��G�/��EMR��l��z� L       split_indices[$l#L       {                         
   
      
                               	                     	   
                  	                            
                                                 	         
                                                                                                                                                                                                                                                L       
split_type[$U#L       {                                                                                                                   L       sum_hessian[$d#L       {F�` F+� E�� F� Dd  E*� EXp Fh D�@ C�  C�  D�  D=@ Bd  ET� E�x EZ� C�� D�` CԀ Bd  C�� B�  D�� C�  D@ C   B   A�  E"� DH  E,  E� C}  EJ� C�  Bd  B(  D�  Cˀ A�  ?�  B`  C=  C&  B�  @@  D�  A0  C�� B�  D� Bh  A�  B�  A�  A�  A0  @�  D�  D�� D� C5  E� D� D�� D<@ B�  C  D=� Ep C  C+  A�  B  A�  A�  C�  D�  C�  A  @   A�  B  A�  B�  B�  @�  C!  A   Bx  B�  D�� @@  A   C$  C?  B�  Ap  C]  C�  B(  A�  A`  AP  A�  B�  A�  @�  A  @�  @@  A   @�  @   D(� DS� C� D� C�� Cr  B  C  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       123L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       mA�R�C'=�s�C�N����FL� ƕ�C9�#Fݤ�F����|�F�/�����"5�3��AFǜF<>HlFR�G-���h�Ƙo�ER6��t�G��G�ě��B%Ǝ��ǩ�_CW���.��?�FޝG� H�ԊG���M҇E�H GZ��F�s;�D���E�3��ʮ�F:�F���ǥ�#G�G~FH�dDu�G�2EmA`Ʃ�o�1>�G��F��J����B��D���dđ1f�x��F5�NŪ��śiCF*��(�'F���F��G�@7D���Gp�ҙ�C�[u�{��E��E���F����H�gF��@���I�ŧR�ƅ]E�7���uI�7��c�.F�H���F��tĐO��	'���F�r�FU�Ţ�E��'����F�g���]FJE=Ɓ��F�F��G�sƮ��Śe��8���J��L       
categories[$l#L       "                            	   
                                     
                                         L       categories_nodes[$l#L             	            "   (   6L       categories_segments[$L#L                                                                !L       categories_sizes[$L#L                                                               L       default_left[$U#L       m                                                                                                 L       idi1L       left_children[$l#L       m               	                     ����               !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _��������   a   c   e   g   i   k����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       mP�\�P�f�Q&1�Qb�AQ��Q-��QnGaP�oR$�TPn�>Q3��Q$ �    P�T=Qb^Q	�_Q��Q�OlQ�4PLp�P_6P�	Pv[�Q~ P�hBP6�PN3Q���Q��FPƟ�Q��Q��Q6��P��P�@�Q���Q�P�P�XN�KTNL��P�0�P�N�P�YCPϗ�PcM�OJG�P�`P@�        PY��P��Q-7$Pd�O�7�NCk                                                                                                                                                                                                                 L       parents[$l#L       m���                                                           	   	   
   
                                                                                                                                   !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   3   3   4   4   5   5   6   6   7   7   8   8L       right_children[$l#L       m               
                     ����                "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `��������   b   d   f   h   j   l����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       mA<z�?��>cS�?̬?���?��FA   @kC�      @�  >49X���?���@�  @��?p�`B�G�D��    >P�`@�F@[�   >�t�A�=q   A�  Bb�\?��HB���>�R>��B8     D�` >�r�@@  @�
=BD�   B�33@?+@G�P@@  D�� =�`B=Ƨ�?��TDu�G�2?�t�@�  B�
=   >���C  B��D���dđ1f�x��F5�NŪ��śiCF*��(�'F���F��G�@7D���Gp�ҙ�C�[u�{��E��E���F����H�gF��@���I�ŧR�ƅ]E�7���uI�7��c�.F�H���F��tĐO��	'���F�r�FU�Ţ�E��'����F�g���]FJE=Ɓ��F�F��G�sƮ��Śe��8���J��L       split_indices[$l#L       m         	      
         
              
                	                                       	      	                                                 	   
                       	                                                                                                                                                                                                                   L       
split_type[$U#L       m                                                                                                     L       sum_hessian[$d#L       mF�` F�� CK  F�T C݀ Bp  C  F�� B�  B  C�  Bh  @   B�  BX  F}� Cl  A   B�  A�  A   CW  CA  AP  B4  @@  B�  B  A�  FyD C�� B�  C  @�  @@  A�  B  A  A�  @�  @�  B�  B�  B�  B�  @�  @�  A�  A�  ?�  @   BL  B  A�  @�  A@  A  Fxp BT  Cw  B(  A`  B�  A�  B�  @@  @�  ?�  @   A�  A   @�  B   ?�  A   A0  @�  ?�  @�  @   @@  Bx  A�  B  B�  B�  A  B@  B,  ?�  @�  @   @�  @�  A0  A  A�  B<  @�  B   @@  A�  ?�  @�  @@  @   A   A   ?�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       109L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       qA�j��=��C��CK  �\�F���C���E"�g�i(F�P7���AF���ǜ��7��Cɕ��=,7E_�eƆ��F��2EC��G�p� ��F��Ǥ�G
����%F�x��$���v<G,F�C�{dǹ\`EР/Īt!FLX������d�'@ Fa���7�LF��H(���@h�L>.�m�9G�eVƇ�MF?.�����Ff��G�ȖFzz�7F�F_��`XDũ���51CG������	B��8F��̯�[(F��<Ŵ�E_��!�5E��Ƭf�ō��EɅp�hN�D�)D�.gĀ��ƹh�E�9F���Ŗ�eEb73Gr��Eڐ��_�7�5�GE���Ű�+��iĹ�gF�څF[�Ƃ7����`�Fq5ŇU�G��F(0{E����؛ND��M��0F��<Ť;Ǉ���XE�]G�y�����Ŀ�y��RLD�ѾED������L       
categories[$l#L       E             	                          	                                               	   
                                                                       	   
                                      	   
            L       categories_nodes[$l#L                                         !   %   )   ,   .   0   1   2   7L       categories_segments[$L#L                                                  	                                          #       %       &       )       ,       .       6       7L       categories_sizes[$L#L                                                                                                                                            L       default_left[$U#L       q                                                                                     L       idi2L       left_children[$l#L       q               	                                    !   #   %   '   )   +   -   /   1����   3   5   7   9   ;   =   ?   A   C   E   G   I����   K   M   O   Q   S   U   W   Y����   [   ]   _��������   a   c   e   g   i   k   m   o����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       qP�s�Qh��P�ÐQ6�`R�lQdg�P�/tQY��P���RdXQ�xQ���Q^^Q}P�QU�vQTAFQH@eP��O��JQ��;R�"R�Q��mPݤ�Qs:�    NmɚQ��R��R
�vP���P�;�Pf} Q(�RQ���P�}&P��L���    QrS�Q�N�QX��P&�Q�%�RiPP��Q@t    N���P���Q�V        P��7Q5�jP��QrDR.[~P���Pؘ�Q� �                                                                                                                                                                                                                L       parents[$l#L       q���                                                           	   	   
   
                                                                                                                                   !   !   "   "   #   #   $   $   %   %   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   0   0   1   1   2   2   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <L       right_children[$l#L       q               
                                     "   $   &   (   *   ,   .   0   2����   4   6   8   :   <   >   @   B   D   F   H   J����   L   N   P   R   T   V   X   Z����   \   ^   `��������   b   d   f   h   j   l   n   p����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       q=���B���=��T   =P�`B�  =0 �@   D�� =49XA   =�PA  B��{=L��?��/   D�  @�  B���   >�I�   D� A�  ��%            B�           ?;d?�A      Fa��>���B���   D�@ >�P   =���   F?.�         Fzz�7F�?�n�B=�H   @?\)>�M�=e`B@�  A`  �̯�[(F��<Ŵ�E_��!�5E��Ƭf�ō��EɅp�hN�D�)D�.gĀ��ƹh�E�9F���Ŗ�eEb73Gr��Eڐ��_�7�5�GE���Ű�+��iĹ�gF�څF[�Ƃ7����`�Fq5ŇU�G��F(0{E����؛ND��M��0F��<Ť;Ǉ���XE�]G�y�����Ŀ�y��RLD�ѾED������L       split_indices[$l#L       q                                                                                                                   
              	                                                              	                                                                                                                                                                                                                         L       
split_type[$U#L       q                                                                                              L       sum_hessian[$d#L       qF�` D٠ Fq� D�� CĀ B�  Fpd D�� C8  B�  C�� B�  @�  C  Fn  A�  D�� C0  A   B�  A�  C�� B  @�  B�  @@  @   B�  A�  A�  Fm� A0  A   D<  CÀ B�  BL  @@  @�  A�  B\  A   @�  C  B�  Ap  A�  ?�  @�  B8  A�  ?�  ?�  B�  A�  Ap  @�  A`  Ap  Fh4 C�  @�  @�  @@  @�  C�  C�  C�  A0  B�  A�  B  A@  ?�  @   A�  A   A�  A�  @   A   @�  @@  B�  B�  Bx  B8  @@  A@  @�  A@  ?�  @@  A�  Ap  A   A   B�  A�  A   A@  ?�  A`  @�  @   A  @�  @@  A@  FR� D�  C�  @�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       113L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       qAc�CI��ŏ^~E���*��U��FXCǫ��E�h��+�C�������a��s�\G[����F��-�F��eD��>�>d�)"GƈC#xFFd@�ƊEkǸ����.~FX�Ɗ�G����84Fs$GuC��:�QG'lFv���q�7D��f���2G~ĸ_F-D���E���G币E` �ͳ��0��>��ǡ<��ۅG�CẈ�3��H4F)e�F����CRE����Q��F�qh��-��;��OGU �E�Uő�F���ƸH��]��56FLŶ6�#s9Gs�E�J����F���D�8Fup�CLʜ�u��'�RF"��E�zZG=t0���F�(ċn��zI��8@F�p�z�K�E�M��Ķ���!��EԐ�E�k�G!��E�Ծł������i5��3F_��F���G��F'Nz�R
B�G!��zbL       
categories[$l#L       	                               L       categories_nodes[$l#L          	                4L       categories_segments[$L#L                                                  L       categories_sizes[$L#L                                                 L       default_left[$U#L       q                                                                                                   L       idi3L       left_children[$l#L       q               	                              ��������      !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c   e   g   i   k   m����   o������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       qP]a�P��cQ�nQ��-Q��Q���Qq�L40 Q�/�Q���Q��>Q�I�Q�>Q6^R �        Q���Q�� Q�iQ���Q|,�Q
xMQ{�:QͶOP��P�2�P��P�LRL�rQOQN��Q�߈Q��RCQ@�P���QrxGQ¢�Q��vQ���Q�ԼQ�Q%)�P�)Q[ʓQj�PO���N"R0O��Po�
Q�I�P��\Q�,�Pw[�R�x�P�a�    P�%G                                                                                                                                                                                                                        L       parents[$l#L       q���                                                           	   	   
   
                                                                                                                             !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   :   :L       right_children[$l#L       q               
                              ��������       "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d   f   h   j   l   n����   p������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       qA"{=��>�j=��=�j>�z�@@  B�  >�-   =��?�w?��   ?�����F��-�B|ff>�r�   B��3@�  =���?yXBY33>�Q�>\(�D�� A,��   >j~�B\��   B�  =��=��
?�B|ffAp  >�>�oB��{A�  >��@   @��P>uB5\)@�  D�@ @�  B�33   B�  D�� B�B�B���F��E}  E����Q��F�qh��-��;��OGU �E�Uő�F���ƸH��]��56FLŶ6�#s9Gs�E�J����F���D�8Fup�CLʜ�u��'�RF"��E�zZG=t0���F�(ċn��zI��8@F�p�z�K�E�M��Ķ���!��EԐ�E�k�G!��E�Ծł������i5��3F_��F���G��F'Nz�R
B�G!��zbL       split_indices[$l#L       q            
                                                            
                                                       	         
         	                                                                                                                                                                                                                                                             L       
split_type[$U#L       q                                                                                                           L       sum_hessian[$d#L       qF�` F� D(@ D:@ Fv� C�  C�� A0  D7� DT@ FiT C�  B   CD  B�  A   ?�  C  D� B�  D>� Bx  Fh\ B�  C�� A�  A�  B�  B�  A�  B@  B�  BP  D  B|  A�  Bt  D'� B�  B  A�  C�  Fc� B�  @�  C  B�  A0  @�  @�  A�  B  B�  B  B\  A@  A�  @   B8  B�  Ap  BD  @@  D @ @�  @�  Bd  Ap  A0  B  A�  D� B�  B�  @�  A@  A�  A�  @�  C�  B  F8� E,P Bl  B  @   @@  B�  A�  B  B�  @   A  @�  ?�  @�  ?�  A   A   A�  @�  A�  B  B  @@  BH  @�  A  @@  A@  @�  B,  @@  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       113L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       A���B+3D��YE9X����su�E���E�V3�k�]D��G�x�XC6pƀ��E����c�U��*�F$���kG��婕�-YEǭ�ƍSi�K����ZE��JG(�[ƤJ�EԈFGa��Ņ��b�Š��F1��E�:TG y�F��KǱ��(�ǲo�ǘ�D�\E���Ӎ�F/����=�ŵېDT/�F�ŉ&E��G4G��C��nE5W�XHEeF���F3ֹH>��CXƢ�?*;ǈ#��Ƕ[�'nFu���oE��EH�S�p��F�iE�o�F�@�Ō ?��$Fj�E<���D��'�/����]�XAC�)6�Qz�D���FV�wFp'��HߠF�u�ă�Fx���"Ǻ�	;��N�uF&��ì�E�ؽ�0�yƂX|đqhD|��F]$�G�"�F$�TG �tƛ�MF�
?Ō(=E=S�i�Ŷ
vƘG7D_zpF�o�F#o�ö�XƨpHFHE	Gw@�F#s���"�F�aƞ�vD��E�4ƱͲ�{Sŋ�L       
categories[$l#L       G                             	   
               	   
                                   	   
                                                                 	   
               	                                   	   
            L       categories_nodes[$l#L                                  &   +   /   9   :L       categories_segments[$L#L                                                                %       &       '       4       8       9L       categories_sizes[$L#L                     
                                                                             L       default_left[$U#L                                                                                                                   L       idi4L       left_children[$l#L                      	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c   e   g   i   k   m   o   q   s   u   w   y   {   }����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       P\��Q"��Q�(�Q`��Q]֜Q�:�Q�
�Q�7:Q]��QK��Q<��Q���Q���Q�
�Q#�bQ=�Q�kQ���Q^UQ+�QBQ�1�Q9�Q���Q���Q9N�Q��0Q��RS9�P�@P�*,QUʒQO� R#��Q�7�P��aQc`LQL�Q*��P�<\Qh�QI�>QWC5Q�L�Q��FQa��Q�x�Qh��Q�BvQ6VR*�WQ(+�PNu}Pω�Q�VlQ{٨Q� 
Q�t!Pd�P��-P;[�O�TPP;�                                                                                                                                                                                                                                                                L       parents[$l#L       ���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <   =   =   >   >L       right_children[$l#L                      
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d   f   h   j   l   n   p   r   t   v   x   z   |   ~����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       A�  >C��>aG�      >�33   >z�H   @@  >^5?>8Q�   ?&ff>�V?ŁB���>��B���?\)B�ff@9��@�D� >�X      >��yB�=q   >��B���?�~�B���>�33>\(�>�Z>�1   A   A   B�  @      <�9X@��
>��   D�� >�p�D�` @�  @   B|  B�33@^��>�S�      ?C��>�o>.{>ix��'nFu���oE��EH�S�p��F�iE�o�F�@�Ō ?��$Fj�E<���D��'�/����]�XAC�)6�Qz�D���FV�wFp'��HߠF�u�ă�Fx���"Ǻ�	;��N�uF&��ì�E�ؽ�0�yƂX|đqhD|��F]$�G�"�F$�TG �tƛ�MF�
?Ō(=E=S�i�Ŷ
vƘG7D_zpF�o�F#o�ö�XƨpHFHE	Gw@�F#s���"�F�aƞ�vD��E�4ƱͲ�{Sŋ�L       split_indices[$l#L                                           
               
                                      	                      
                                     
          	                     	          
   	                                                                                                                                                                                                                                                                      L       
split_type[$U#L                                                                                                                         L       sum_hessian[$d#L       F�` Ft E� E� E� E�@ E
� E
 C+  E"� E�  E�` C�  D�� C<  D�� D�` A�  C  D�� D�� Cq  E�� EJ� D�  A�  C�  D�� B  C  Bh  D\� Ck  Dz@ B�  @�  A�  C  @�  @�  D�  D�@ B0  B�  C,  E5� D� C�  E,� D�� Bl  A0  AP  B�  CT  D�  C�  A�  A   B�  A0  A`  B0  DS  B  B�  C  Dn� B<  A�  B�  @   @�  Ap  @@  B�  B  @@  @�  @�  @@  De� C�  D�� B  @�  B  A  Bp  A  C#  D�@ D�� B�  D�` C�  C  A�  E+0 D�� A�  ?�  Bh  A   ?�  @   A0  B�  A�  C  B�  D�� A�  C_  C  @�  A�  @�  ?�  B�  A�  A   @@  ?�  AP  A0  B  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       127L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       {A�TLDX֐���ă�mE�VXĭ[F��E���Or0F/��ļ�TB��dŴ��F%>�G�o=D�[�F���ż�2E:��Fj��ƀ��GU�&�+��aF2��F�k�����E�G��z�2��H�VƏnPE$��G,���	�{��OƝ!�F�����F��|Dץ�������H6�������>E����C�ܡD�Z)G��G��B��R��G�Ɖ�D0�>G%��H4l�ú'3G�ƭ��H/��E�PU�a^�ō� E���C���G��F$�"�/��F@��E���ĹG&�9�<��-~D7#F�S�FM7`���F+Ed��ŹUPE��g�s��Sa���f�T��F �G�Y�F����	�!�Vĳ�0�\Y�D��ĄdR�`��Db�P�v;��&iEw�F;�q��AG���Fz*}ľ�F�X��?��EDz\�s=�Ɩ$,Fp �T�_GxO�Fr4�FLTŒ�?Fx��@y4Gd�F.�7F*���L       
categories[$l#L       \                    	               
               
                               	   
                                                 	   
                                            	   
                                     	   
                                                 	   
            L       categories_nodes[$l#L                    	         $   &   '   -   /   7   9   :   ;   =   >L       categories_segments[$L#L                                                                 !       "       .       /       1       =       K       M       N       [L       categories_sizes[$L#L                                                                                                                              L       default_left[$U#L       {                                                                                                  L       idi5L       left_children[$l#L       {               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c   e   g   i   k   m   o����   q   s   u����   w   y������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       {Pbc�Qg!SQ]�Q/��R �sQ; �Q��QdDQj�lRPQQ�aqQ(`Q��QT�FQ�~�Q3r[Q0
�Q�{Q�~�Q���P���R(��Qx]lQ�Q���Q��Q��QV�Q��P��^Q)��Qd��QE��P�:\PC��Q+�tQ���R4zQ��9Q�U R�UP���P��Q��lQP�nQ��QC�Q�Q0Qj#�Q�պQ��Q)�Q��vRc�Qw/m    OP|�O()�Oբ    P� Ob'o                                                                                                                                                                                                                                                L       parents[$l#L       {���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   9   9   :   :   ;   ;   =   =   >   >L       right_children[$l#L       {               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d   f   h   j   l   n   p����   r   t   v����   x   z������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       {   D�  A      ?�r�   >�D?i�^? Ĝ   D�@ B�  @   E}  ?�
@@     B�  @'�@�z�   ?(1'@��D�@ ?�\)D�� ?t9X@<��>�@��?�o<�h@�  D� B�  =o   @        @陚?�?�P@E�>      =�   D�� >!��@�  >�S�@�  ?
~�B�     G%��         ƭ��      �a^�ō� E���C���G��F$�"�/��F@��E���ĹG&�9�<��-~D7#F�S�FM7`���F+Ed��ŹUPE��g�s��Sa���f�T��F �G�Y�F����	�!�Vĳ�0�\Y�D��ĄdR�`��Db�P�v;��&iEw�F;�q��AG���Fz*}ľ�F�X��?��EDz\�s=�Ɩ$,Fp �T�_GxO�Fr4�FLTŒ�?Fx��@y4Gd�F.�7F*���L       split_indices[$l#L       {                       	   	                                            
                           
                                  
               	          	                                                                                                                                                                                                                                                                                               L       
split_type[$U#L       {                                                                                                          L       sum_hessian[$d#L       {F�` FD E�� E�h EV@ E�� C  E` Edp D�  D� E�P D�` B�  A`  E� B�  E� D�� D�� C9  A�  D� E�� C�� C  Dߠ B�  @�  @�  A  B�  E	� B<  B   E  C�  C  Dq  Do� C̀ B�  B�  A@  A�  D:  D�� C�  E�� Ck  B�  B(  B�  D@ D@  B�  @   @@  @�  @@  @   @�  @   ?�  B�  C6  D�� @�  B,  B  @�  B�  Ep B�  C8  B�  B   B  Dg� C�  D� C?  CZ  B   B  B�  Ap  @�  @�  @@  A�  B�  D  A�  D�  C�  Bp  E*  E� B�  C  B�  @@  ?�  B$  B�  @�  D@ C�  D.� B�  A�  B�  @   ?�  ?�  @@  @   ?�  @�  ?�  ?�  ?�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       123L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       B�&D�D�� ĥ�\
E�*�B{�DB8D�R����FYǒŬXE��o��e`��sD�����F�2D�8�ߡ�F	r�G5�FVI��Sy�C��F�v�A۝ƒi�Ǆ)Ė_@��E�7&����D%��F7BG�B�F��qőrIG{���Ej~G�tG�����D�;TG�j��WW�`�GKyq�)R�FXGZZq�  �D�hE����Åu����*�Fj����ΐ(D%XM��Fv�F��!�vDF����u�CH�OFbv��$GL�/F
���ANN���F$�x�2��F�>5�"��ƃi�Eυ�]Fr[2���	G
�F8qƈ�F!p�G��E|��WGw>E��Ɨ��Š��E��G	�]D�G�Ŏ�nD*�&E^F��E��G hD��jŮ���pF;�F���쮧�����Ca���Ɖ�x�o	��c�ĦY�Fa�*�Blg��.�&zF3��E.˯�$^�Z��Ɛi:F�`�ElҳL       
categories[$l#L       7                      
                                                  	                          
                     	                                  	   
               L       categories_nodes[$l#L       	                         /   2L       categories_segments[$L#L       	               
                                   "       (       6L       categories_sizes[$L#L       	       
                     
                                   L       default_left[$U#L                                                                                                                     L       idi6L       left_children[$l#L                      	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c   e   g   i   k   m   o   q   s   u   w   y   {   }����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       Ps.;Qz�Q?Qb��Q�$hRLpQQ3MQ��xR+U#R(�Q�aeQ��Q��:Q��6QEg�QP�1Q�`Qw��RfQ�q�R
R�RR|Q-��Q��QG�Q��Q{��P���Q�O�Q��Q<Q<Q�^R[:nQ`Q+Qtd&Q��WRӖQ���Q�ΎQ�z�Q���Qz�Qq0�Q-$Q~[�Q<�AQ)ߦQ�lR2�VQ���QZؕQ�� Q��PNјP�*@P���P��(Q�i�Qk,Q�H,Q��                                                                                                                                                                                                                                                                L       parents[$l#L       ���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <   =   =   >   >L       right_children[$l#L                      
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d   f   h   j   l   n   p   r   t   v   x   z   |   ~����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       >XbD�  >��yB���>�1   >S��Bq33   >�ȴ>��yB{��B~=q>Y�A�  <���Bd  =�\)   >��   >�bN>��#=�\)@���>z�HD�  B�     >�`B>�$�      >��H?(��>���?�E�>aG�>��wD�� B$  >R�@��@   =Ƨ�B�R?���   =��wB�     A�  B�  =�
=D�  =�9X@�  >��9B=�HA�  >��?��>���F��!�vDF����u�CH�OFbv��$GL�/F
���ANN���F$�x�2��F�>5�"��ƃi�Eυ�]Fr[2���	G
�F8qƈ�F!p�G��E|��WGw>E��Ɨ��Š��E��G	�]D�G�Ŏ�nD*�&E^F��E��G hD��jŮ���pF;�F���쮧�����Ca���Ɖ�x�o	��c�ĦY�Fa�*�Blg��.�&zF3��E.˯�$^�Z��Ɛi:F�`�ElҳL       split_indices[$l#L          	      	                          
                                  
   
   
      	                
                          
                  	                                                 	      
                                                                                                                                                                                                                                                                L       
split_type[$U#L                                                                                                                             L       sum_hessian[$d#L       F�` E�p F5 E�p D�  E�( E�� EJ� Di  Dm� C�  D�� E,  B�  E� E:� C~  D � C�� DM@ C  C  C�  D�@ Cɀ D�� D:@ A�  BD  E�� D�  B�  E50 Cc  A�  C5  C�  A�  C�  D/� B�  B�  B,  B�  A�  B�  C�  A�  D�@ C�� Bx  D,  D�� C  D� A�  @�  B  Ap  C&  E�P C�  D)� AP  B�  E� D&  C/  BP  A`  AP  C   BT  CԀ B  A  A�  B�  C  C;  D � B�  A�  B   BX  A�  A�  A�  B�  @�  AP  A   Bh  C  B�  @�  A   C2  D\  C�  @�  B,  A�  C�  C�  D�` B  B�  B�  A�  D@ A   A0  @@  @�  A�  A@  A@  @@  C  A�  D8@ E�H C�  A�  B  D   L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       127L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       sA��p÷FZEP��!��� 4|E��~�k!�C����OE��c�G3��FO���^e��H���śE�ޣ@>'D]����)F��ƫVGij���&��q�F�3�ƥ�0Gk�Ǒ�YF2�F���Ķ�QF_�dƁَE�d���<��{��E���FT�_�Gø�C��Ɔ��ǱipG&� GBl�D�k�ٿ�E����CF�F��ƅ�z���mGx4tF���<��ŕ�T
kF 6�G��,������H2EF_qE薾�yE-�8q�EP�F7�fD��.�����\�F�=gM��1Fw�D"�X5E`}E٭�ŝ�?G"qFE�E2���j����E3in�|��/S�F\���J�MFj������C?�FR�G�L�)B�E��aF�>�����E7A��6y$�-�F�T����ũ~�{��Â_�Ŷ�4G���Iƪ�j��Ea��ŃR�E����Ӻ�L       
categories[$l#L       M                           
               	                                	   
                                                            	   
                                        	   
                                              	   
         L       categories_nodes[$l#L                	                  #   '   /   0   1   7   9   =L       categories_segments[$L#L                                                                       "       #       $       /       0       >       A       BL       categories_sizes[$L#L                                   	                                                                                    L       default_left[$U#L       s                                                                                              L       idi7L       left_children[$l#L       s               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W������������   Y   [   ]   _   a   c����   e   g����   i����   k   m   o   q����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       sPYr�Pډ\Q:��P��Q�	nQ�TgQ6f�P� �Q��Qv�Px�TQ��~Q��,PՑQ& �Q�FhP� _QY��Q��|Q�2�Q���P��HN��|Q�T�Q��.Ql�|Q�@�O���O$kNRo�Q"��Q���Qc5�QZ~>P���Q�XQ3,Q$mQY��PR��Q5��QIQ0�|Oy�            Q6P�vxQ~��R:LQ�)P((�    P﮲NG@    MF��    Q�:
PJ��Q�z�Q��p                                                                                                                                                                                                                L       parents[$l#L       s���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   /   /   0   0   1   1   2   2   3   3   4   4   6   6   7   7   9   9   ;   ;   <   <   =   =   >   >L       right_children[$l#L       s               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X������������   Z   \   ^   `   b   d����   f   h����   j����   l   n   p   r����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       s?�?G�>ٙ�      ?�9X>���=��`BVff   @33D�@ B�  ?.�D� >��=ě�>"��   ?;d@�  >�V   ?��B=�HB�(�B�ff>{�m      @��   >�5?=�%@+S�   >_;d?��@@     B�  >���D�` @ĜGBl�D�k�ٿ�         ?!%@ĜA33Gx4t?;d   �ŕ   F 6�@���>�~�   @�=qE薾�yE-�8q�EP�F7�fD��.�����\�F�=gM��1Fw�D"�X5E`}E٭�ŝ�?G"qFE�E2���j����E3in�|��/S�F\���J�MFj������C?�FR�G�L�)B�E��aF�>�����E7A��6y$�-�F�T����ũ~�{��Â_�Ŷ�4G���Iƪ�j��Ea��ŃR�E����Ӻ�L       split_indices[$l#L       s                     
   
                                                              
                                                  
                             
          	                                                                                                                                                                                                                                             L       
split_type[$U#L       s                                                                                                   L       sum_hessian[$d#L       sF�` Fb� E(� F]� C�� Df� D�@ FA D� C�� A�  D;� C,  A�  D�  C�  F9� D� DO� BH  C_  A�  @�  C:  D  C  A`  AP  @�  B�  DҠ C�� B�  D8@ F.$ C(  DU� CW  D  A   B(  CR  AP  Ap  ?�  @   @   B�  Bp  CU  C�� C  @�  @   A@  A  @�  @   @@  A�  BL  D?  Df@ Cl  C  BP  B,  BD  D,  F-� A   B@  B�  B|  DE� AP  CJ  B  D� @�  @�  B   @   C  B\  @�  @�  A`  ?�  A�  B�  B`  @�  @@  CR  C�  B�  B�  B$  @@  @   @�  @�  @   @�  ?�  ?�  A�  @�  @   BD  CL  D  C�  D @ L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       115L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       {A��nÎ)�E#���{�������F/*bÚ�yF>hFV���p����FX��F�џ�-�k���fƮ��F�=�ƈ�WĐ��Gt`AǾ�
E�]�D�7���Gv?�b�MHD�&F��@D݀��u�����FE�X%��u�Jx�G@���ƀ}��(F�j��8C;Gl�G���D�@ �(��ԣG��Aƈ$��_'FGU0�vJ�Ǚ�%H�G�>F1g�CHf�E��)�F3�4G`T���Gi� �f%n��BI���E;.�my�-�E����V���@lFK�rG��C~�7���D�9FƱ7��'�6F8�'��4Ń�G9"{D�trł��G!�ņ	�Fg�GEÐh�~ǚE�%��=	F���E_�3�)AZFA���i����F�ªEV������ޡ���e��n Gs�F,K��+ʿF=h��f�E�Q����Ņ?�E�MgG��`E@6G!��Ť��G��Œz�E�4&F�2EMG��c;QF�o�L       
categories[$l#L       3                      	                                     	   
                                                                     	   
                         L       categories_nodes[$l#L       
                  %   +   -   0   1L       categories_segments[$L#L       
               	                                   !       "       /       0L       categories_sizes[$L#L       
       	              	                                                 L       default_left[$U#L       {                                                                                                          L       idi8L       left_children[$l#L       {               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c   e   g   i   k   m   o����   q   s   u   w����   y������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       {PMKQ�"�Q��Q!�R+$ Q�~�Q��0Q��dQ�tQ-�"R��RB�*R Rw��Q��
P���QԽ�RQ��Q�СQ���QŠQHĠQ�+Q�o�R7��Q���R��Qw$�Q���QV�
Qg8ZQ%�Q�� Q�"%Q٨bR$:&Q�r�Q��P�LQ9hAQȪQ�JO���P"�Q=`P!¼P���Q�,xQ���RlR7��Q*�Qky�Q���Q���Q(    R	�xR=cQQ^-�P���    P�R�                                                                                                                                                                                                                                                L       parents[$l#L       {���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   9   9   :   :   ;   ;   <   <   >   >L       right_children[$l#L       {               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d   f   h   j   l   n   p����   r   t   v   x����   z������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       {B���B�B�D�� B�  D�@ >�+   B�=q?Z��A�  @'�?�G�>�ƨ=8Q�A  B�        ?b>��      @�ff?Qhs@�  >��D�  B�  A   A   @   B���D�� >n��>�\)?D�D�     >���?A%>���>���@�     =�t�   @�  A�      >�B�(�>��>��j@��
>J��)�@�  >��/Ap  B�(��f%n?JBI���E;.�my�-�E����V���@lFK�rG��C~�7���D�9FƱ7��'�6F8�'��4Ń�G9"{D�trł��G!�ņ	�Fg�GEÐh�~ǚE�%��=	F���E_�3�)AZFA���i����F�ªEV������ޡ���e��n Gs�F,K��+ʿF=h��f�E�Q����Ņ?�E�MgG��`E@6G!��Ť��G��Œz�E�4&F�2EMG��c;QF�o�L       split_indices[$l#L       {                            
                                                      
                        	                                                               
                	             
                                                                                                                                                                                                                                                L       
split_type[$U#L       {                                                                                                                 L       sum_hessian[$d#L       {F�` Fp< D�  Fn< C   D�� D$� Fi� C�  B|  B�  DI@ C�� C�  C�� Ff� C?  C=  B�  BD  A`  B(  A�  D� Cr  C   Ci  @�  C�� C{  A�  FY� DM� B�  B�  C  Bd  B�  A�  A�  A�  A   @�  @�  B  @�  A�  C�  B�  C-  B�  @�  B�  C;  B8  @�  ?�  C�  B4  Cl  Ap  @   A�  FFT D�@ D<� B�  B  B�  A�  B`  C  @   B0  AP  A�  B  @�  A�  @�  A�  @�  A�  @   @�  @�  ?�  @�  @   @   B  @@  @   AP  @�  C� A  A�  BL  C  A�  A�  B<  @�  @@  A0  B�  A�  C   A�  A�  ?�  @�  C�  A   A�  A�  C	  B�  A   @�  Ap  ?�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       123L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       kA��LūX�C#u+FL���m�g��bWD��G��QF$�m!��!���@G>&�FCJC�G?|�Fc�+F�iaƇk�"ւ�EYGoƅN�Dm��žk-G�\FÄfE��HG�6�ǀٲCB��FIM��D�F:_�G�Q���3���D�o{��=�x���GXk�Ƒl��/D���Dd�G��ŋϯǺ�bG<0E2��Fu��E��CHv�F��U�@� G�7����h��)F��yB��F�d|E/�G3�wEM��E��Y�L�E���Jݭ�P�w�%EF�K����yƇ�tǁ33�>�F�HEo$N�v@�E��oƊt��ȡ�*Ć�E�IFT��G@�š]�ÈQIE9g��.�~FW��Ť�E���'��͇SF9:�F	J�AW�E���G%i��	'�*��D�e~F�:��Y)�BX��L       
categories[$l#L       !               
                                            	   
                                         L       categories_nodes[$l#L                         $   &   .   4   7   9L       categories_segments[$L#L                                    	                                                  L       categories_sizes[$L#L                                                                                    L       default_left[$U#L       k                                                                                            L       idi9L       left_children[$l#L       k               	                              ����      !   #   %   '   )   +   -   /   1   3   5   7   9   ;��������   =   ?   A   C   E   G   I����   K   M   O   Q   S   U   W   Y������������   [   ]   _   a   c   e����   g   i����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       kPB�MQ��PRU�Qw��Q�L.Q+�Q��mPģtQ)șQ<�Q��nQAiP�g�R�FQ"�{    Oj=�QD��Q3PXP�V�P�Z�Q�aQ%��Q�iR6}.P]�O���Q��Q�X�P��P�@�        P�� Q\�pQ7�0P�0P�P�P|�N��     P�WP(��Q�Q�eQ<ÛP��Qa�Q��            P 3Q��*Q�ePI��Q�� N    Q@�Q�p                                                                                                                                                                                        L       parents[$l#L       k���                                                           	   	   
   
                                                                                                                     !   !   "   "   #   #   $   $   %   %   &   &   '   '   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   4   4   5   5   6   6   7   7   8   8   9   9   ;   ;   <   <L       right_children[$l#L       k               
                              ����       "   $   &   (   *   ,   .   0   2   4   6   8   :   <��������   >   @   B   D   F   H   J����   L   N   P   R   T   V   X   Z������������   \   ^   `   b   d   f����   h   j����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       k=t�   >�R>o>�b?�>,1@�     >u>��@XQ�=� �D�� D�` G?|�   B�  B��@�  @�  @�  ?8Q�?�+BD     @   B  =�
=   D�� FIM��D�=�C�? ĜD��    >���   Bv{���<uD�` =�hB�  ?��
   @��R>F��G<0E2��Fu��   >�I�@@     B7��   ��)Bd  D�@ F�d|E/�G3�wEM��E��Y�L�E���Jݭ�P�w�%EF�K����yƇ�tǁ33�>�F�HEo$N�v@�E��oƊt��ȡ�*Ć�E�IFT��G@�š]�ÈQIE9g��.�~FW��Ť�E���'��͇SF9:�F	J�AW�E���G%i��	'�*��D�e~F�:��Y)�BX��L       split_indices[$l#L       k          	            	                  
                                                                                 	                    
                                                                                                                                                                                                                                                 L       
split_type[$U#L       k                                                                                                L       sum_hessian[$d#L       kF�` Cр F� C  C�� EL� FS @�  C  B  Cq  EK� A�  D � FK @@  @   B�  B4  A�  @�  B  CL  D�  D�  @@  A`  C�  B  A  FJ� ?�  ?�  B�  A0  B(  @@  A�  A   @@  @   A�  A  B0  C   D�@ @�  D�@ A�  @   ?�  @�  A  C�� B�  A  A�  @�  @�  B  FJ\ @@  B�  @�  @�  A�  A�  ?�  @   A�  @   @   A   ?�  @   @   A�  @�  @�  A   B  C  @   D�� D;  @�  @   C�  D�  A   Ap  @@  @�  C�  B�  A   B�  @�  @�  A   A�  @   @@  A�  A   A�  FJ L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       107L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       A��|Ĩ��D��EԄ��(ED�>��(R��!��Fzx�PBE�PpFrD
e��D�D�:F�|�Վ~GP�{F-.X�GZƄ0F�8cE�AF��q�#���8��EɃŔK����~�pb'E�aG������G�.�}%)�MG�ŜFdk�����3�[F�>�Eޔ��/G�-�ĵ�u��J�E� �Db�G++�ƫ��F�wBD��z�{	GR��E�s�<pE�M�[	P�M��F�\��`F-o��X�2{1F��E�ƭ�E�t7Ɗ 3��`���|�F+�g�Y�G
s�E���ż�E����"W�Ɗ����ѣņ��GK�E�o�<ȵF��;�7��FS�����F�؝�2x�E)��F�{��O��Ea-�����E���y��Fi�2ƅ����:E{D�F����D����F�ġg-G8d�G,A�FD� WF�M�"%��n�F���W�Q�q���-3�ELq�?���b�F=�NE�c��|��C�w�E�|�Ɠ�|�QL       
categories[$l#L       P                               	   
                              	                               	   
                  	                                                  	   
                                       	                                  	   
L       categories_nodes[$l#L                                      '   3L       categories_segments[$L#L                                           $       '       .       ;       ?       E       GL       categories_sizes[$L#L                            	                                                        	L       default_left[$U#L                                                                                                                     L       idi:L       left_children[$l#L                      	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c   e   g   i   k   m   o   q   s   u   w   y   {   }����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       PJo;QF
P��Q��^Qf�Q\j Q6<Qm	8Qk�.Ql|xQ.�0Rf�;QL�Q�{QXQ�FzQJ �Q1L�QF8Q�E!Q���Q�>hQg&�RA�XQ�FQ(8Q��jQ&�.Q#�4QgJ�Q^�Q{q�QhP
Q���Q�PP��"Qb�Q=�ePm�QOQ�LQQ�H�Rt�Q� PM�$Q�޻Qb,�Q��R��QT>�R��8Q%��Q�Q�Qh��Q8T�QQ=T�P�P��PQ�0eQe�QpJP,~1                                                                                                                                                                                                                                                                L       parents[$l#L       ���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <   =   =   >   >L       right_children[$l#L                      
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d   f   h   j   l   n   p   r   t   v   x   z   |   ~����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L          >|�?��T>o?�u   ?�X      ?�l�D�@ @J?-   @�  =�hs@�  B6ff@�G�@M�T   >��>/�D�� @��@��   >�33BZ        B@  >7K�B(  >M��@�  B���>8Q�>��   =�Q�B�G�A  B8��D�� ?�$�?�>���?X��?��F@fv�   BL  >ۥ�?�ĜB�ff?hs@��R?�
=?�Z>=p�BP  D�  �2{1F��E�ƭ�E�t7Ɗ 3��`���|�F+�g�Y�G
s�E���ż�E����"W�Ɗ����ѣņ��GK�E�o�<ȵF��;�7��FS�����F�؝�2x�E)��F�{��O��Ea-�����E���y��Fi�2ƅ����:E{D�F����D����F�ġg-G8d�G,A�FD� WF�M�"%��n�F���W�Q�q���-3�ELq�?���b�F=�NE�c��|��C�w�E�|�Ɠ�|�QL       split_indices[$l#L                
      
                  
         	                                                                       	                                  
                         
   
                                                                                                                                                                                                                                                                                        L       
split_type[$U#L                                                                                                                           L       sum_hessian[$d#L       F�` E�� F<� D@ E�P F� E@ C9  C�  E}� D  DJ  F� D"@ D�` B�  B�  B  C�� Ei� C�  Bl  C� C� C�� E�� D�  D� B�  DS� D@ B<  B  B�  A�  A  A�  C�� A�  Ed  B�  B�  CK  A�  B  Bp  C̀ CK  C~  Cz  B�  E�  E� B   Dx  C�  CN  B|  B`  Cr  D  C�  B�  A�  A�  A�  Ap  B4  A�  Ap  A@  @�  @�  A`  A�  B  Cy  A   A@  EL� C�  A   B�  B�  A�  C6  A�  @�  A�  @�  A�  A  BL  C�� B�  B�  B�  Cp  A`  CT  B  B<  BX  EL` E'� E` @@  @�  A�  Du@ A0  C�� A�  B`  C  A�  B<  BD  @�  C9  Bd  B�  D � CO  C�� @@  B�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       127L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       SA�}`�W�B�)F��ƹ�C!�xŹF��5Ft��8�F�|Cf�F�и�Pk�\@x�
�FM�AF����GG�GY�9��C'~���g�G�?i�{����� �n�AŰ�G�'D���a�F(|Sæ� Ef�.�p�-G`XvţRU� ��E"��B�'�F0Fua��=G	0�E���шG%V��۝4��tƳC���1s��V�E+Gm�E`�D�%������ƨ2�F��'E���DJi4�E����XTEQՀ@�f�E��>F@��6wƔ9��b_D�Z�}����g�<�rEj��F�p�Mcg�"ؚD0�Q�$)�FBĵ��L       
categories[$l#L       %               	                                                               	   
                                  L       categories_nodes[$l#L          	   
                   #   $   (   ,   2   4L       categories_segments[$L#L                             
                                                         !       "       #L       categories_sizes[$L#L                                                                                                  L       default_left[$U#L       S                                                                 L       idi;L       left_children[$l#L       S               	      ����                        ����      !   #   %   '   )   +   -   /   1   3   5������������   7����   9   ;   =����   ?   A   C����   E����   G   I   K������������   M   O   Q������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       SP+��Pћ�PWO��xP�QjP�giP���    O��P�erPL
Pu�P��O���Q=��M��v    OJFP��O�*ROFϖPp�TP���P�WNP� �Kp�(OVb0PE��PUtP            ME��    PG��M�6@M��    N�^P�C*QEOh    P���    K�^M��`N��(            MS��O�5PE��                                                                                                                        L       parents[$l#L       S���                                                     	   	   
   
                                                                                                                 "   "   #   #   $   $   &   &   '   '   (   (   *   *   ,   ,   -   -   .   .   2   2   3   3   4   4L       right_children[$l#L       S               
      ����                        ����       "   $   &   (   *   ,   .   0   2   4   6������������   8����   :   <   >����   @   B   D����   F����   H   J   L������������   N   P   R������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       S=m�hB"  ?�p�?�ff>P�`@��>�+F��5B��      @7L?I��=�Q�@�C�   FM�AB0�\=#�
A�  B9��?�9XBff   BK��   ?a��@�F   D���a�F(|S   Ef�.@@        � ��@�  @�F   Fua�D�� G	0�   B\)B�33�۝4��tƳC�   BNG�   Gm�E`�D�%������ƨ2�F��'E���DJi4�E����XTEQՀ@�f�E��>F@��6wƔ9��b_D�Z�}����g�<�rEj��F�p�Mcg�"ؚD0�Q�$)�FBĵ��L       split_indices[$l#L       S         	                                                     	                                                                                                                                                                                                                                             L       
split_type[$U#L       S                                                                      L       sum_hessian[$d#L       SF�` Bl  F�� A   BD  F�� C�  @@  @�  B  Ap  F�� A�  A@  C�  @�  @   @�  A�  @�  A  F�~ A�  @�  A   @   A   C}  @�  ?�  @�  @@  @@  @�  A�  @�  @   @@  @�  F�| C  @   A�  @�  @   @�  @�  ?�  ?�  @�  @�  A�  Cc  @@  @   @   ?�  @�  A�  @@  ?�  ?�  ?�  ?�  @�  F�$ B0  B�  Bx  A0  A0  ?�  ?�  ?�  @�  @   @   @   @   @�  A�  A   CY  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       83L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       wA�Ѿ��:C��R��u�`%mF�8B�K�F�o�I�?F:��ƤPF�j~�K3�D�H��∯F�|�ŊȔ�V>��)|E�|�GI���m^R�p��E�6G)�+�C�D�0�ųy�Eba�E�B�C�F�$�H,TC<,�aV��ފ^�;��ȨǎF)��'y<E��MF�	��UѮ�����D�v�FY��PтǄq~GC<	ƈ��ǰ�kFc�pa��hŚ�]�|P�E���E]d�G%6��f��\�&E�˙Fl��G��f�W�4�i�E�����R
F��L�5�;�+�&��C��r��ő��'E���%i�ƒ�oŌ�����F݄J�#�v^��O�"�Y��F�d��i�wF��F�ƯG�ƾ���4F8vEG�Ǝ�&DD���!�� ��F��5�E{���XE������f�'�2ݥD�q�E��F�%�C��PĲ<�F�#.�OZ4Eڧ���e�FE�GL       
categories[$l#L                                     	   
                                                            	          L       categories_nodes[$l#L       
                      (   1   5   8L       categories_segments[$L#L       
                                                                       L       categories_sizes[$L#L       
                                                               	       L       default_left[$U#L       w                                                                                                  L       idi<L       left_children[$l#L       w               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G����   I   K   M   O��������   Q   S   U   W   Y   [   ]   _   a   c   e   g����   i   k   m   o   q   s   u��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       wPEdQHP�P�̻Qw��QF͛QWMOP]�^Q���Q f�Pv��QR$�Q�c<P��Q*��P�gQ�y�QN��Q�VQ��Pe�wN� Q,�Q��Q_�Qk�P��Q[�QfTQ$��Qe3�P��Q4�Q0�hQ5�:Q�_�OZ�    Q�FP<��P2�O��0        QD�Q��|QY�PX4�Q	�P₼OS��Q[��P�tRO"� P��-P�މ    QC+Q8;�QM�bQQ׫Q��3Pщ�Q��|                                                                                                                                                                                                                                L       parents[$l#L       w���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   %   %   &   &   '   '   (   (   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   8   8   9   9   :   :   ;   ;   <   <   =   =   >   >L       right_children[$l#L       w               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H����   J   L   N   P��������   R   T   V   X   Z   \   ^   `   b   d   f   h����   j   l   n   p   r   t   v��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       w=\D�  =��   B{   > Ĝ>��j<�h?�x�A�  @@  @@  >%=��T?D�B�
=   ?j=q?E�T>=p�>G�?C��BVff=D��   ?ƨ<D��=�>��A�        >�$�=���A0  �;�=�9X?ٙ�>p��   E��MF�	�=���=Ƨ�?�/B�  B  =�h   A0  D�� D�     @@  ��h   @�  B�  =�B4z�C  BP  E�˙Fl��G��f�W�4�i�E�����R
F��L�5�;�+�&��C��r��ő��'E���%i�ƒ�oŌ�����F݄J�#�v^��O�"�Y��F�d��i�wF��F�ƯG�ƾ���4F8vEG�Ǝ�&DD���!�� ��F��5�E{���XE������f�'�2ݥD�q�E��F�%�C��PĲ<�F�#.�OZ4Eڧ���e�FE�GL       split_indices[$l#L       w                               
            	   	                
         
             
                                         
                  	   
         	                                                                                                                                                                                                                                                                            L       
split_type[$U#L       w                                                                                                             L       sum_hessian[$d#L       wF�` E� FgP E� C�� C�  Fa� C� DȀ Bt  Cr  C,  CD  EZ� F*� C�� C`  Ap  DƠ BT  A   CU  A�  B�  B�  A�  C*  D� E2� C�  F$D C�� @   CO  A�  AP  @   D�� @�  B@  @�  @   @�  A�  C<  A�  A@  B�  Ap  @�  B�  A�  @�  B�  B�  @@  D� B�  E,0 C�� B4  F!� C  C[  B0  ?�  ?�  B�  B�  AP  @�  A  @�  D� D~  @�  @@  A�  A�  @   @@  Ap  A   @�  C6  A0  @�  A0  ?�  A�  B4  @@  A@  @@  ?�  B�  A   @�  Ap  @   @@  Bx  B  A�  BL  B|  D  A�  B�  E$p B�  A�  C�� A�  A�  F! B@  C  A�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       119L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       w@�PD�]Ø+E+p�H��DX���@C��F�=F�r��W?ĀzlEk��V�՟ME~$����E,�F�U���=�G�gǒz�Ʃ5�EԻ��F
 ïN�F!J�t� E�U�q��C�E�F��ǬJw���U�CF�Gb��FW߆G��#w�E�u������˻���HE�r�Gw�a�ۭ,��-OF.*��=U�G9Qčw;Eӈ'G�n���#F�F]̟ŧV?�Y����Db����_Fh\�\N�����DF� �6��F�l�ő1�E���WHF�L�E�\�FD��G0E���E�$Qƀf����E�FV��J�F�|iŋw�EK+��J�D�r�Fխ��ŉ�Ģ%mDMͶă��E�V�t�V�B���F���C���[�Eh���Z0�E�gG9iæ!2���F����c�F'aE�F��3�$EbuXŰu�Klx�-~L       
categories[$l#L       %                       	                                                                              	   
             L       categories_nodes[$l#L       	                       $   &   /L       categories_segments[$L#L       	                             	                                   $L       categories_sizes[$L#L       	                                                               L       default_left[$U#L       w                                                                                                        L       idi=L       left_children[$l#L       w               	                                    !   #   %����   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O����   Q   S   U   W   Y   [   ]   _   a   c   e   g   i   k   m   o   q   s   u����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       wPX@Pמ�P��yP�a�Q��oQ'��Q\QH7[Q�2�Q!.^P��QD�Qh{P��FQִ�Qm.�QX�QF?hQl8"    Q�%�P���PO�<Q�3NQ��Qr��QDs`Q���P� �Q"eZQ�)�Q��tR ��P�Q5O�QUԤQ��dQQt�Qp��P�|lP��    O���P�)P�*�QKX�Q �Q*sQ4�Q��rP���Q��Q']�Qu�;P�H�QC��Q��|Q��P���Q��}Q',`                                                                                                                                                                                                                                        L       parents[$l#L       w���                                                           	   	   
   
                                                                                                                                   !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <L       right_children[$l#L       w               
                                     "   $   &����   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P����   R   T   V   X   Z   \   ^   `   b   d   f   h   j   l   n   p   r   t   v����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       w   ?��   ?�{   D�  A�  >��
D�� >vȴ?���=�7L?�r�=��   B���@   >5?}@b��=�?��HB  BHA�  >Y�   D�@ ?f��@�  @�  B�  B�\)   @��=���=\)   ?H��   D�� @�K�E�u�@   >�@IG�D�` @@     ?*~�B$ff?�p�@�  B�aHB�  @�  A0  >   >hr�=��D�@ >5?}Db����_Fh\�\N�����DF� �6��F�l�ő1�E���WHF�L�E�\�FD��G0E���E�$Qƀf����E�FV��J�F�|iŋw�EK+��J�D�r�Fխ��ŉ�Ģ%mDMͶă��E�V�t�V�B���F���C���[�Eh���Z0�E�gG9iæ!2���F����c�F'aE�F��3�$EbuXŰu�Klx�-~L       split_indices[$l#L       w      	                            	                                	                                           	                                            
                                                                                                                                                                                                                                                                            L       
split_type[$U#L       w                                                                                                              L       sum_hessian[$d#L       wF�` E  Fg@ E0 B�  F� E�� D�� D)@ B   B�  E�h E:� E�8 D�� D�� C�  D� C  @   A�  A  B�  D� E�� D�� D�@ C^  E�H C�  D � Dg  CP  A   C�  C  C�� B8  B�  A@  A�  @   @�  B  B@  D� A�  D�` Eu� D�  C  A�  Dʀ CX  @�  E�� Cu  Cy  CQ  D@ A   DV  B�  B�  B�  @�  @�  A�  C�  @@  C  C  CU  A�  A�  A0  B�  A   @�  A`  @�  ?�  @�  @   B  A�  A�  C�� C'  A   A�  D)� C�  D�@ E� C~  Dn� B�  Ap  A�  A@  D�@ C�  CD  A�  @   @�  E�8 B�  B�  C  Bt  C<  A�  C:  B�  D@ @�  @�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       119L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       s@�ŵ��B���Ey��Տ�Ff-�B������Gp��~F���G0H�����^ƘB�΃G3fsť�*� ��G��mż���|WG�5��o�H9mFm���C�UF��ƥI�GV�Eӣ8�A� G����/�Eɼ*ƅ�IG�|ǆ��GO�#G_��Ƽ�OGh�nƏ��Ǭ��Gw��F0@��\�G�"Gb#GK��G8�6�Z���qX�ƚ,gFV's�ej �'��Ee���=U�G��EBhGKD�ŒN+Cx�����gF�1ET��{5�ƃ [Ea�E 4�48F�Y�œr�Ş����%LF��HF+�F�:���F��<ĵ�MF�2�0P,�^����8!ZF���E��=���D�}F�'3�C��F���F2�A���Ƣ#��}��F?��(�Dǔg�K��k%�E��0F|H��aFֺE�h'� �Fm�YĻ��F��g�����+E�4pBBCL       
categories[$l#L       .                  	                                      	   
                                                       	   
                           L       categories_nodes[$l#L                            #   (   6   7   =L       categories_segments[$L#L                                    	                     )       *       +       ,       -L       categories_sizes[$L#L                                                                                    L       default_left[$U#L       s                                                                                             L       idi>L       left_children[$l#L       s               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I����   K   M   O   Q   S   U   W��������   Y����   [   ]   _   a����   c   e   g����   i   k   m   o   q����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       sP0�QY TPI�Q"�Qd�>Q��GPAv�P�Q�l�Q_��P�_�Q��;P��jP�OJPc&�P�x�P�NXP��.P��$Q�Q+v4P<M��(P��HP݀
O���O:<�P��P��Qr^P��'P�,�O�SQ��Q�O���P"��    Pa��Pw`LO���Pu Q
ߘO�l�N��        O2`    P��FP��zN��O�j    Mo�P\X�Pb�X    Na7�Q�Q��Q���P�(�                                                                                                                                                                                                                L       parents[$l#L       s���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   $   $   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   /   /   1   1   2   2   3   3   4   4   6   6   7   7   8   8   :   :   ;   ;   <   <   =   =   >   >L       right_children[$l#L       s               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J����   L   N   P   R   T   V   X��������   Z����   \   ^   `   b����   d   f   h����   j   l   n   p   r����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       s=49X   =D��B�B�>Õ�   =P�`D�  >ؓu?�T?Vȴ   ?ŁB4  =��>�A�>��yB�33   >���   D�� @ۅBM\)@��@-   ?��D�� B���=�jA�  B�
=��B7��   >oGO�#@   =���   ?�z�>p��B  Bq33�\�G�"B  GK��@�  D�  D�  >�-FV's      @��R�=U�A   D�` D��    =�����gF�1ET��{5�ƃ [Ea�E 4�48F�Y�œr�Ş����%LF��HF+�F�:���F��<ĵ�MF�2�0P,�^����8!ZF���E��=���D�}F�'3�C��F���F2�A���Ƣ#��}��F?��(�Dǔg�K��k%�E��0F|H��aFֺE�h'� �Fm�YĻ��F��g�����+E�4pBBCL       split_indices[$l#L       s               	             
      	      
                                                                  
          
                                                                                                                                                                                                                                                                                                      L       
split_type[$U#L       s                                                                                                        L       sum_hessian[$d#L       sF�` C�� F�� Cz  B�  Bx  F�: Ca  A�  B�  A�  B  A�  Bx  F�� A@  CU  A  A�  A�  B(  A`  @�  A  A�  A�  @�  Bd  @�  C�� F� A   @�  B�  B�  @@  @�  @   A`  A�  @�  Ap  A�  @�  @�  @@  @   @�  @�  A`  A�  AP  @�  @   @   A�  A�  ?�  @�  C�� A�  DX� Fr� @   @�  @   @   A   B�  B  B�  @   ?�  @@  @@  @�  A  ?�  A�  @�  ?�  @�  A0  A`  AP  ?�  @�  @�  @   ?�  @@  @�  A   @�  A@  A   @@  @   @�  ?�  ?�  A�  @@  @�  A�  @@  ?�  C�  Ap  A`  A`  B�  DB� B�  Fq� L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       115L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       uA��9ĖAD	��Ek��?��E�|��c~�E΋��7�ż\aEG0~E�RkǠ�j�W��BF�ƫ��c��GR���E3# ��ϛF�[�E���F��MČ����E�k��I��Y%�F�&�F>L�đ�nF�����SY��8��Ű�#G�T!ƕ@Ť�^F�,/�gG���FW�G�t�(�\F"p�i-�FM�G�m�F~�!�jF����~ISD�Y�G����Y�G�=đ��E:nCG-�Ɓ�8E���DȡcE�Q��E�ō��Ƙz�l=Fl�yEb���q��ŔP�F�]F�1�����w��$_�2|�C��yEU8Fx��R����V(��'�Dv�(�U�E���F$�jGL|XE���,��E���D���XE���E;�G%i:G,�ZD�u��2�m�(��FVf� �F�K�Ć��[A��n�}ń���l���D����4W�F��t��S�F�}9L       
categories[$l#L       ;                              	                                     	   
                  	   
                                                                         
                L       categories_nodes[$l#L       	                   $   '   7   9L       categories_segments[$L#L       	                                           "       *       .       :L       categories_sizes[$L#L       	              	                     	                            L       default_left[$U#L       u                                                                                                        L       idi?L       left_children[$l#L       u               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A����   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c����   e��������   g   i   k����   m   o   q   s������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       uP&�pP�N�Q9�,Q��FQk��Q�V'QyQ��Q���QB�&Q�,=QS�Q���Qdg�Q6�=Q,D2P���Q�=�Qxn_Qh�vQ7QaQ���Qp"Q�`PZ�WO��P�URQB8P�I$Q�7Q?rQCa1    P�QQ��ZQTb�P�P�(QYJ�Q��Q>qoP��^Q�!Q���Q��bQuT�Q�5�Q/J Qy��Q���    M�        P��Py��Q*e�    Q��Q�|�Q�JXQ)                                                                                                                                                                                                                        L       parents[$l#L       u���                                                           	   	   
   
                                                                                                                                         "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   4   4   7   7   8   8   9   9   ;   ;   <   <   =   =   >   >L       right_children[$l#L       u               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B����   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d����   f��������   h   j   l����   n   p   r   t������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       u> ĜD�` >C��B�  By33@�  ?\)>���B�  >�~�@�
=>�S�   B5\)B�  ?��   >�G�=P�`>���>��9B$  B�� D�� B�B�   A�  ?\j>�A�A�  @�        F���@@  >���   >�+>ۥ�   >^5?BH?
=q>ݲ->&�yB�  @#ƨ@�  A   A�  ?���F~�!?������~IS   B     G�=D�` B&ff>��>x��E���DȡcE�Q��E�ō��Ƙz�l=Fl�yEb���q��ŔP�F�]F�1�����w��$_�2|�C��yEU8Fx��R����V(��'�Dv�(�U�E���F$�jGL|XE���,��E���D���XE���E;�G%i:G,�ZD�u��2�m�(��FVf� �F�K�Ć��[A��n�}ń���l���D����4W�F��t��S�F�}9L       split_indices[$l#L       u                                    	                    	      
   
                                                 	                          
                     
                                      
   	                                                                                                                                                                                                                        L       
split_type[$U#L       u                                                                                                            L       sum_hessian[$d#L       uF�` E�@ F:� D�  EUp D�� F"� D�� C�  E� D�  D�@ A0  CG  F� D�� B�  C�  B(  D� D � DU� Cr  D�� C;  @�  @�  B�  B�  F� C  Df� C�� @   B�  C�� B�  A�  A�  Cր D�� B�  Cɀ D%� CA  C   B�  D;@ D� C&  A�  @   @�  @@  @   B�  @�  B�  ?�  E�H E0 B�  Bd  C�  C�� B�  C�  B�  Ap  C�� A�  A�  B�  A�  ?�  A�  @   C  C�� DN� D	@ B�  B  A�  C�� Cs  Cр B8  C  B�  @�  B�  B  CS  D� C�� B�  C#  @@  AP  A   @@  ?�  AP  Bl  @�  @   B�  B`  C[  E�p D� Dـ A�  BX  BX  @@  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       117L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       OA�h2��XQF�H�ÿ��D�<�F����r�����Ś�*E�)����RéjgG 	ź���wg�Ò=8G (D[�qƢ"�GJ�E����X�E(E�GDD�I�D䬢ą�7���G�j�w��F�SD���R1D�уG�%IEї�Ƌ�EE���ƙ�G�D���G6��Fr1 @09�EJ.1�gEKŁ��E ���.DGl4JE���F7b�8F�l�D�dĄ�Gk"N�D��)�F%�$ŶY�GpV�F�S��xlES6�F���ȑ�E��E�+���$���7˙GC�FE�P����Fm�D��4E�����D�L       
categories[$l#L       %                                                	   
                            
                         	   
         L       categories_nodes[$l#L                      !   (L       categories_segments[$L#L                                                  L       categories_sizes[$L#L                                                 L       default_left[$U#L       O                                                                    L       idi@L       left_children[$l#L       O               	                  ����   ��������               !   #   %   '   )����   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       OPCY:PC�O��.P�8�P�}TO2�L���Q�k,Q��=QT�Q
�9    N���        P�K�R�w�Q�k�R/TQ��}Q'�Q��Qh�3N���    Q]��QkrQ��R���Q�Q�-�Q�(R��P�P�Qy��Q?0�P���Q�W�QZ7�Qz"Q��N�3�Nl�                                                                                                                                                L       parents[$l#L       O���                                                           	   	   
   
                                                                                                                 !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *L       right_children[$l#L       O               
                  ����   ��������                "   $   &   (   *����   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       OA�  ?�   B�  >ٙ�=�j   B�     >ȴ9?=p�éjgB�  ź���wg�>� �?9X>�p�?�?�/?��D�@ ?D�>D��D�I�B�ffB�  @z�   >uD�� ?�  >gl�   @@  D�@ >$�/>ݲ-Be33>��T   >Q�B8��@09�EJ.1�gEKŁ��E ���.DGl4JE���F7b�8F�l�D�dĄ�Gk"N�D��)�F%�$ŶY�GpV�F�S��xlES6�F���ȑ�E��E�+���$���7˙GC�FE�P����Fm�D��4E�����D�L       split_indices[$l#L       O                                
                     
   
   	      	                                         
             	   	             	                                                                                                                                                   L       
split_type[$U#L       O                                                                         L       sum_hessian[$d#L       OF�` F�< A�  FbH E(� A�  @   FV$ DB@ Df� D�@ @   A`  ?�  ?�  FU B�  D  CQ  B�  DU� D� D�� A@  @   Ed0 F B  B   C�  B�  B�  B�  B   A�  DB� B�  C�� C�  B`  D�� A  @@  E=� D  F� Cb  A�  AP  A�  A�  Bd  CԀ A�  B`  B�  @   A   B�  Ap  A�  @@  A�  C;  D  @   B�  B�  C/  C2  B�  ?�  B\  C@  Dq� A   ?�  @   ?�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       79L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       yA��cC����2C{��F�6Ficp�0�����WC�FE0�G
���a�GG�ī��ƃz�����E�ZF%�>C��,G�����E�"��G�K��_a����G"�%�27���Ɔ�@�82C���ƚC���V�G��jĉl��i�GM�E�K��F�S>Hi��~pE4HEF��'����Gʚ�ţIKE#�U�` |E8�'G�;���|FR%kű��E�eƬ��G��N�u&����/ƚ,GG}����!H@�������F�G�%5Ű�kE��Ű��E};DE���GM EHO"C|VA�g�.עFMh[���GI��F��=�����x��F�^�PU�8dF�Ԥ�^R�?9gGO�qP�F�a#ƚ-$�`�pFF�y��]���E�z��9c�F�u��+\��tM�',�F�.'��h�D9�ŏ�lė� E$�%LE��dD���G�L"Ūް��Y#�ŞF,Y�D�^��b�hE��G#+xL       
categories[$l#L       ,                        	                                               	   
                                              	   
             L       categories_nodes[$l#L                         &   (   .L       categories_segments[$L#L                                                                +L       categories_sizes[$L#L                                                               L       default_left[$U#L       y                                                                                                              L       idiAL       left_children[$l#L       y               	                                    !   #   %   '   )   +   -   /����   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c   e   g   i   k   m   o   q   s   u   w������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       yPT_P�u�Q@Y�P��aQO��Q�x(Qe�Q���P���Q�&Q��AQ��Qcs\Q�nQ�(=Q}� Q�n�Q�K�P�4Q$��Qt| Q�niQ�W�P�B�    Q���Q�Q4�Qc�:QȝQ���P�J�P[g�Q���Qb<�Q#�5R��Q)7�Q,<oO��N�� P�Q"f�QVؽP�HQ}��QQ��QwNP�>%P�� QYT�O!��P*��Q���Q>r�Q3�Q���Qt��QQkçQaF�                                                                                                                                                                                                                                                L       parents[$l#L       y���                                                           	   	   
   
                                                                                                                                   !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <L       right_children[$l#L       y               
                                     "   $   &   (   *   ,   .   0����   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d   f   h   j   l   n   p   r   t   v   x������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       yA�  A�     ?�G�>�l�>Kƨ>�{   ?��RD�@ D�� >�n�?��?�$�>�ff      >�A�>E��Bn  =49X   >Ƨ�A  ���@@  D�� >���?���@@  B���>�33D� A�  >dZBX  Bk��? A�   @�     @D�� B��{D�� A     Bx  >��wB�  @�  B�=qB  ?��R?��\?�7BJ�>e`B>�ĜBH@�  ���!H@�������F�G�%5Ű�kE��Ű��E};DE���GM EHO"C|VA�g�.עFMh[���GI��F��=�����x��F�^�PU�8dF�Ԥ�^R�?9gGO�qP�F�a#ƚ-$�`�pFF�y��]���E�z��9c�F�u��+\��tM�',�F�.'��h�D9�ŏ�lė� E$�%LE��dD���G�L"Ūް��Y#�ŞF,Y�D�^��b�hE��G#+xL       split_indices[$l#L       y                      	               	   
      
                           	                   
                                                             	                                                                                                                                                                                                                                                                                    L       
split_type[$U#L       y                                                                                                                 L       sum_hessian[$d#L       yF�` FZ� EH� FT� C�� C,  E> C�  FO  C�� Bx  B�  B�  E,P C�  C  C]  C_  FK� A0  C�  A�  B  B�  @   B�  A   E$ C  C  C  C  A   A   CS  C'  B`  E�  F
 @�  @�  A`  C�  A�  @�  A�  A0  B�  @�  B  B@  @@  @�  Db@ D�  B�  @�  B�  B�  B�  BX  B�  B�  @   @�  @�  @@  B�  B�  B�  B�  B  A�  D@ Edp FD D  @�  @   @@  @   @�  @�  B8  Cf  A�  @�  @�  ?�  A�  @�  @�  @�  BL  A�  @�  @@  A�  A0  B0  @�  ?�  @   @   @@  C�  Cπ D<� Dq� B�  A�  @�  ?�  A�  B4  B@  A�  BH  B$  BH  @�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       121L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       mA� UDT���s��C��rFh��4�J���iY�Eϗ'F���t�G?���B�DEd<��sD��6�bp�Eo�F�H8G�G�F���E+������q���;F�x�E���Qm�E��tD�)��ݍ�s�QG�
G֚EV@�G?Z�F;1ƐyGܦ�ǞF�F�5G��yĕ�`ƺ,0�2.1Cp��Ǖ�F�.���l�h8�F��{F$�Cs�E5����D�FP����C2t�E&��F���11�D�����Gi*F2gD����$��Ey��F���E��eħT�E�<Z�1�'G'O D�K�F#0���|F�[�E���G{b��-�*E�S2�p�ůC�E�T�E�[ŗ[��sE���F]V6ƌQƣ������J�����G!g�7uTEgFq�=D��H�l}E�`�æ��F6&���|De/�F*�;F�B�YL       
categories[$l#L       6                     	                                  	   
               	            	                                                                 	   
             L       categories_nodes[$l#L       
         	   
         "   %   )   2L       categories_segments[$L#L       
               
                                   !       &       '       5L       categories_sizes[$L#L       
       
       
                                                        L       default_left[$U#L       m                                                                                              L       idiBL       left_children[$l#L       m               	                  ����                  !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?����   A   C   E   G   I   K   M   O   Q����   S   U   W   Y   [   ]   _   a   c   e   g   i   k����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       mPS��Q�,FQ�JP�HoQ�k�Q�
0Q,	~Q�wQ"SuQ��P�\E    Q���Q�ЯQ`ΞQ#�Q�& P��	P��Q��bQ��mP��PP��aQ,s$Q`�Qa�QW��Q��4Q�JpQD]�QO;�Q	��O��    P��Pg��O��O��Q���P�-�Q{�RQj��P�+'    Oη�Q��P�><Q&Q)��P��DQY�Q�	�QgP�Q��eR�Q�@tQ�                                                                                                                                                                                                                L       parents[$l#L       m���                                                           	   	   
   
                                                                                                                                   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8L       right_children[$l#L       m               
                  ����                   "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @����   B   D   F   H   J   L   N   P   R����   T   V   X   Z   \   ^   `   b   d   f   h   j   l����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       mB\  BX  Ba��@X �   <�t�   @�p�BP        G?��   >\)?b   @�  D�� >�ƨ@�  ?L��?s33=ě�B�  >$�D�  B���D�  @Co@@  >&�yB�R>�+G֚   D�� @      @��H>�\)>���   @�  ƺ,0?*~�?Ͼw>�o@�  >�I�B��{   A33D�� >k�<���?˅@�{C2t�E&��F���11�D�����Gi*F2gD����$��Ey��F���E��eħT�E�<Z�1�'G'O D�K�F#0���|F�[�E���G{b��-�*E�S2�p�ůC�E�T�E�[ŗ[��sE���F]V6ƌQƣ������J�����G!g�7uTEgFq�=D��H�l}E�`�æ��F6&���|De/�F*�;F�B�YL       split_indices[$l#L       m                                                  	                               
                                                                 	      	                     
      
                                                                                                                                                                                                                   L       
split_type[$U#L       m                                                                                                   L       sum_hessian[$d#L       mF�` F� E�0 F0 C�  D  E�P F� D3� CC  C  @   D� E@ E�� E� E� D  B�  A�  C'  B�  B  C�  Cp  BD  E0 E� DD� E�� D� E� @�  ?�  D� B  B,  @�  A�  @�  C!  @�  B�  @�  A�  C�� @�  A�  C^  B  A@  Dl@ D�@ D�� E/` D   C�� E�� Dg� B   D
� DC� D�  @@  @   C�� C  A   A�  A�  A�  @   @�  A�  @�  ?�  @�  A�  C  ?�  @�  A�  B�  A�  @�  C`  B�  @�  @   Ap  @@  A�  CC  A�  @�  @   A   D_� BH  Dk� C�� C�� D�@ B�  E*� C�� C  A�  C  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       109L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       yB%m��ȳC����$e��FE���Ì��E��.�}�IEÅ��G�F7L�Q�C���ŏkE�j��HY�����@�F7���G�D����&��G4�E��G�4�ŀ�����F&��E����
_�G-�D��ƽ�O�PȌƉ���q��GA�Ţ7�E~�GI�F�S,ż�EWZ�-�Ɔ�4F�T�G�@Gִ�EF} F�g����G1&�ſ�hFd�DE���"�E G;igF�C��u�ŐJO��fF_�Y�����E��O�w>.Fd��%�l�'���cB���F́%�еE�K,ŸjRE���RӬG /E�mC�^#F��K�_��4�E8GR�C�E�~ŉ�1�)4��GAeEpFT ŅcG�S<FO�F���D8L�F�2ER����-Zƺ���HF7k����D��ŋ�Q���b��F��FJYF�)�EBFF��-��!Ƣ���j�E��z�6k�F^��L       
categories[$l#L       3                     	   
                     	                     
                                                                           	   
            L       categories_nodes[$l#L             	               -   .L       categories_segments[$L#L                      	                                          %L       categories_sizes[$L#L              	       	                                          L       default_left[$U#L       y                                                                                                       L       idiCL       left_children[$l#L       y               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C����   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c��������   e   g   i   k   m   o   q   s   u   w����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       yP0�4P�K�Q�lQ�K�QM�Q�k�P��Q\/QdZBQ3�
Q_u�R	��Qo�,P���Q�rQ9NQU��Q���Q�CQ�gP��6P��[Q㝐Q]�QKP��FP�!�P�EQ�ovQ ��Q���QI��Q f�Q�_    P��Q�"�Q��Q<�Q<�dQ�itP�͏P�'�P��P�rxR�R.��Q��Q�d�QWd�Q�Ѕ        P�n�QguQt�Qi:�Q&�Qf-.Qz��P�,UQ�h�Q�y�                                                                                                                                                                                                                                        L       parents[$l#L       y���                                                           	   	   
   
                                                                                                                                         !   !   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <   =   =   >   >L       right_children[$l#L       y               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D����   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d��������   f   h   j   l   n   p   r   t   v   x����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       y>!��=��w>XbD� >��   A�  >�=��   B[z�?\(�@�  A�        B�  B�  D� B�ff      D�  >�7L@�  A�  ?�/?�/>hr�>�%@�  @E�D�� B^  �PȌ?3��>�l�>ix�>O�D�  @   D�@ B��q?)��=T��      @�  >I�@   >+���G1&�?�>��j>���>E��B�  D�` >gl�>�G�>z�HA   F_�Y�����E��O�w>.Fd��%�l�'���cB���F́%�еE�K,ŸjRE���RӬG /E�mC�^#F��K�_��4�E8GR�C�E�~ŉ�1�)4��GAeEpFT ŅcG�S<FO�F���D8L�F�2ER����-Zƺ���HF7k����D��ŋ�Q���b��F��FJYF�)�EBFF��-��!Ƣ���j�E��z�6k�F^��L       split_indices[$l#L       y   	      	      
          	   	                                                                                              	                                      	              
                  	                                                                                                                                                                                                                                              L       
split_type[$U#L       y                                                                                                                 L       sum_hessian[$d#L       yF�` EY� FVL D2  E-P E F5 C�� CЀ Dg� D�� D�� D8� F� D�� C�  A�  C�  C  D� C�� D�� D)� B�  D�� @�  D7� F  C�  C�� D�� BD  Ce  Ap  @   CT  B8  A@  C  C�  C  A�  C�� Dv  C7  D� C  B�  A@  D�� C0  ?�  @@  D&  B�  E�� Ep C}  B\  C�� A�  D]� C   B0  @�  C,  Bd  A0  @�  C  B�  A�  A�  A   @�  B`  B�  C  C�� A�  B�  A�  A0  C�� A�  C�  D� A�  C'  C~  C�� @�  B�  B�  AP  @�  A   A   D�� A�  C  D%  @�  B  B  E�� D�� C�� D�@ Ct  A  B(  AP  C�� A@  Ap  A  D>@ B�  C  A@  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       121L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       sB��Ė\PD��F��\Įo�D�����6GUC��A1��P-DըDy�F���E�Rv�bܺF���G��M��YyE���ļ� �3���{?�E��3DJs�F� (G�KyEڏ�F���.	�Bm�+�(�LşeG>�BGI�F���j���l��ģǬ�L�53w�ɒ�E���Ɯ4$D��F�F&D��iům	Gx�dCH� HL�3G(s�G���.�lE,��F��Ųg��R�_Em��ū��ƈD)V�E�>�ű�F�^aE� t�- �Ek�ē��D�x�C�9��!5��u2���@�N�VF<.�DqzAF�md�>�f�q�/Eo��*U�~��F'sjC��vEsK�ĀlŰ�E��mG1�Jƪ��D��F��G���E��F�GwF�uE����vh��8�]�9��E��PFA>PEG�g�M1�E�3����Ɲ[�E�F�C/*����M��a� ņ�(FEy���WL       
categories[$l#L       #                          	                   
                         	   
                        	              L       categories_nodes[$l#L       	                      &   9   :L       categories_segments[$L#L       	                                                          !       "L       categories_sizes[$L#L       	                                                               L       default_left[$U#L       s                                                                                                L       idiDL       left_children[$l#L       s               	                                    !   #����   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?������������   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c   e   g   i   k   m   o   q������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       sP&�gP蛼P��P��6P��Q
��P�o,P��lO�VtQ-�Q>�Q�Q�7�Q ��QA��P�NO���O�!#    Q)�
Q��vQ�5�Q�yQ-�VQ��RQ��_QH�vP���P���Pɧ�Q=�O&b�O\�            M�XCQ<��P�ETQQ���Q��Q��]Q��XQڶQ��P��uQ�Y]P}#P��P�,Q!�.Q|��Pa�P���P FgO�`hQ'�P�&WQ�JQ��.                                                                                                                                                                                                                        L       parents[$l#L       s���                                                           	   	   
   
                                                                                                                                   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <L       right_children[$l#L       s               
                                     "   $����   &   (   *   ,   .   0   2   4   6   8   :   <   >   @������������   B   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d   f   h   j   l   n   p   r������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       s   >L��?��>?|�>��D>���B  >�>���@���>8Q�?���         BB�RD�  <�E���@u/@�33=���A@  ?��T   @�     @��D�� @@  ?;"�D�` Bv{GI�F���j��B4z�@j=q   ?E�TA  @ ��>�-@�  ? �?$ZB�ff@@  =0 �B@��D�  @   B�  B�
?.�?xQ�??}      @@  ?L1E�>�ű�F�^aE� t�- �Ek�ē��D�x�C�9��!5��u2���@�N�VF<.�DqzAF�md�>�f�q�/Eo��*U�~��F'sjC��vEsK�ĀlŰ�E��mG1�Jƪ��D��F��G���E��F�GwF�uE����vh��8�]�9��E��PFA>PEG�g�M1�E�3����Ɲ[�E�F�C/*����M��a� ņ�(FEy���WL       split_indices[$l#L       s                        	            	                                       
                                                      
                                                                                                                                                                                                                                                                                       L       
split_type[$U#L       s                                                                                                          L       sum_hessian[$d#L       sF�` E�� F<� A�  E�� F E
� A�  A0  EC� D�  Fl B�  C�  D�� A@  @�  A   @@  E 0 D� DX@ D�� F, B�  A�  B�  C0  B�  D�` D'  @�  @�  @�  @   @�  @�  E� @�  B�  C�� D@ C�  DU  Ck  F` D|� A�  BL  @@  A`  B   Bh  B�  B�  B�  A   DB  D� CӀ Cu  @   @�  @   @�  @   @   D�  D%� @   @@  B  B  C� B0  D@ A�  Cx  B�  C�  C�  B�  C(  F� C�� DY  C  A�  A  @   BD  ?�  @   A  @�  @�  A�  B`  @   B  A�  BL  Bh  Bt  A0  @   @�  B�  D$� Bd  C�  B  C�  B  CS  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       115L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       uB	���~-E�B�����tEp�tƹ;È��E�b�
������ĵ>F#uDFI0Fǃ��C.�ŕ�'F�4���o7Ń�G���E�2�T?�e�Ǆ;fFXH��GR�����E��Ǧ��¸ԻF*��F9�G�] �3��F�\2E'�3Ʋx��u6F�s�G�V��i�Gƹ� G1���/��.u�G�m��
1F-y`ǢrTFE��GU"��P3�F�DOG��3GG���m���CĳF��Ǽq���W��nJ�?g�wƣx�Ey�E���ď�YEd Ň���fڣE^��FC����lċU�F-��dx�D�xEF%`i�bϯE�yF�یG+�D�. �L[�F��F��ū���
�x��G���Fk�Ej��.#�E�� D2L���ŭ��ĝ.�Ft+�EW}��#A��G4F��F�X�E6�gE�tƷ��Ƃ��ŀZ�{�AFk?!�K_��i�D�Z���/ML       
categories[$l#L       >                            	   
                     
                                                                                                              
                           
      L       categories_nodes[$l#L                               !   '   )   /   0   1   4   9L       categories_segments[$L#L                                                                                      !       "       )       7       =L       categories_sizes[$L#L                            	       	                                                                             L       default_left[$U#L       u                                                                                                      L       idiEL       left_children[$l#L       u               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S����   U   W����   Y   [   ]   _   a   c   e��������   g����   i   k   m   o   q   s������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       uP3�Q��Qv�cQ.�Q��~Qg�1R
2qP�ʡQ�6Q���Qz�PQ��Q�y�Q�Q��QuOQ��Q��UQ$�XQ��R+�Q��QU� Qy�zP�u(Q��OQT͊Q�qyQk��PZ�IP�I P^A�Q` �Q\��Q�{�Q��Q�]�QHQ���Q�<Q�y�Q�+�    P��PͮS    QO��Q��QY��MP��P�QtQ�9�Q[�        Q�     Nja�P�a�M�\@O��P���N�/                                                                                                                                                                                                                        L       parents[$l#L       u���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   +   +   ,   ,   .   .   /   /   0   0   1   1   2   2   3   3   4   4   7   7   9   9   :   :   ;   ;   <   <   =   =   >   >L       right_children[$l#L       u               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T����   V   X����   Z   \   ^   `   b   d   f��������   h����   j   l   n   p   r   t������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       uB���B�\A�B�     >��T   B���   B�  D�� >���A  >k�@   @�     @@  >��?�D�@ D�  >���>&�y   B�  ?�$�?A%      ?4��<��
=� �   =���>�P@�  ?�>���   @�     �i�G>aG�@�  �/�@            A  >7K�   GU"��P3�>n�G��3   >��#D�� @�  >vȴB�  �nJ�?g�wƣx�Ey�E���ď�YEd Ň���fڣE^��FC����lċU�F-��dx�D�xEF%`i�bϯE�yF�یG+�D�. �L[�F��F��ū���
�x��G���Fk�Ej��.#�E�� D2L���ŭ��ĝ.�Ft+�EW}��#A��G4F��F�X�E6�gE�tƷ��Ƃ��ŀZ�{�AFk?!�K_��i�D�Z���/ML       split_indices[$l#L       u                                                                                     
   	               
                                  	                                                             
                                                                                                                                                                                                                           L       
split_type[$U#L       u                                                                                                      L       sum_hessian[$d#L       uF�` Fp< D�  Fd� D7  D�� B�  FY� D-  D@ B�  Dn@ DC@ BH  B$  FFT D�@ C�  C�  D@ A�  A�  B�  Di� A�  DB  @�  A�  A�  A   A�  FA� C�  C�  Dz� C  C�� C*  B�  D@ B�  Ap  ?�  A�  A0  @�  B�  B  D`� @@  Ap  C  D  @�  ?�  A�  @   @�  A�  @�  @�  A�  @�  B�  F@ A   C�  C  B�  Cn  D?  B  B�  C7  B�  C  A�  B`  B`  B  C�  B�  Ap  A   @�  A`  @�  @�  @�  A   B`  ?�  B  C�  C�  ?�  @   A   @�  Bp  B�  C�  Cb  A@  A@  @�  ?�  @@  Ap  @@  ?�  @@  @@  A   A�  @@  ?�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       117L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       QA݃CF��j�A+k�E���ŇsG��CE�5�.�G�!�Ep�bƏXCyr�B��G0TeEMC�0�	G8@DgGf�E2F�Ƥ�?GR~�0�eE� �CT���9G�8�Fy$���RGA�-ǀ�qF�dG�QF��>�J�F"^sƊ�4�n�Ŕ�F��!�� �F��DDP�8B02�Eڗ�ĸ�ƋoD�))GUGD�D�F�=F���ĘU���F���e+��^�G�/�(��
pgFF�?�x�v�E�?B����t�(�v�� �*��ҮE�1��ɰ���V������ȓû�wF:��ĄGPœ D�H"L       
categories[$l#L       2                               	   
                                    
                                     	   
                     	                        L       categories_nodes[$l#L       	   	   
            "   &   '   )L       categories_segments[$L#L       	                             &       '       -       .       /       1L       categories_sizes[$L#L       	                                                               L       default_left[$U#L       Q                                                                  L       idiFL       left_children[$l#L       Q               	   ����                              ��������   !   #   %   '   )   +   -   /   1   3   5   7   9   ;����   =   ?   A   C   E   G����   I   K   M   O������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       QP%G�PG-�Q\d
P�!QE�Q0�    QϨMQ�ONP~QXQ
�[QA�Q/hP�V�Q�yMP�=�Q�{�        P�i�P�%%P��HP�0�P��P�G�P��hQN&�Q�׌P���P�ܺPFXTQ�DZQl1M    P��P̾OQ`��P��.PlrpO
��    Q{�P�κQ9`�P���                                                                                                                                                L       parents[$l#L       Q���                                                     	   	   
   
                                                                                                                             "   "   #   #   $   $   %   %   &   &   '   '   )   )   *   *   +   +   ,   ,L       right_children[$l#L       Q               
   ����                               ��������   "   $   &   (   *   ,   .   0   2   4   6   8   :   <����   >   @   B   D   F   H����   J   L   N   P������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       Q?��?��FA0  ?�9X<�1@�G��?�%B�ff      D�  @�33@?;d   AP  B�  G8@Dg?�dZBi��@�C�@   @@  @@  @:�\A�  D�     D�  A�     @�  G�Q   Bfff>և+>�+      F�   >�"�?�p�?�;dB02�Eڗ�ĸ�ƋoD�))GUGD�D�F�=F���ĘU���F���e+��^�G�/�(��
pgFF�?�x�v�E�?B����t�(�v�� �*��ҮE�1��ɰ���V������ȓû�wF:��ĄGPœ D�H"L       split_indices[$l#L       Q   	               
                           
                                       
                                                          	   	                                                                                                                                                L       
split_type[$U#L       Q                                                                        L       sum_hessian[$d#L       QF�` F�� D9  Fv� D*@ D8� @   Fr� C�� @@  D)� C5  D@ Fq� BX  C;  B�  @   ?�  A0  D&� C/  @�  CW  C�  Fl� C�� Ap  B  C.  AP  Bd  Ap  @@  A   C�� C�  C#  A@  @@  @@  A�  C9  B�  Cj  Fl$ B(  C�  A�  @�  A  B  @@  @�  C)  @@  A   A�  B  @�  A0  @   @�  C�� A   C   C*  A�  C  @�  A   ?�  @   @�  A�  A�  C  B|  B4  BX  C4  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       81L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       aA�9C�"����Fv��C�iFiG��fF��c�6Ԝ�K�iC�DiE�+OG�g��F`�FD}G���FTSbD��#�kǆz���tE�`C�b�I��F�Yb�k*pG,mī���M�0F�_G!n�G%�G,��F����F��Ɩ��<��E��ƶ�oŖXZFl��ūg���.xCY�VE��3�I���G6$E�A��|GE"Ů���%]qǺǗsFFW�F�>�Ew{�F�z�Dk�ZƲT�E�:�F$�jū�5� D.C�4ř�TƁ'�D�}kF��E����d�A�'uF�zC����v�_E8�ƴ���m����E��-ƃ��Ź��F�D
�NF�2�D��M�u�FŃkF�
��
��F�O��Ÿ���F�Aj�L       
categories[$l#L       ,                            	   
                                  	   
                               
                               	   
   L       categories_nodes[$l#L                   *   ,L       categories_segments[$L#L                                           #L       categories_sizes[$L#L                     
                     	L       default_left[$U#L       a                                                                                           L       idiGL       left_children[$l#L       a               	                                    !   #   %   '����   )   +   -   /   1����   3   5   7��������   9   ;   =   ?   A   C������������   E   G   I   K   M   O   Q   S��������   U   W   Y   [   ]   _����������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       aP"�P��P�_Q	|�P��Q�;�P��QM&�P'wO��P`�9QzQY�fQ.�uQpvNP|5 Q�JP�uO��xN�D    Q�XQ�b5P���Q:�O4�6    Q��Q�?�Q-c�        OO%4P���P��O�:9N⑮Nxi�            Q��JP�Q��?P\alPS�oP'�<P�_>Q��        Q�eQ��Q��mQU-�O�4pP��!                                                                                                                                                                L       parents[$l#L       a���                                                           	   	   
   
                                                                                                                 !   !   "   "   #   #   $   $   %   %   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   3   3   4   4   5   5   6   6   7   7   8   8L       right_children[$l#L       a               
                                     "   $   &   (����   *   ,   .   0   2����   4   6   8��������   :   <   >   @   B   D������������   F   H   J   L   N   P   R   T��������   V   X   Z   \   ^   `����������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       aB   =#�
      D�` ?{A  A0     ?��`D�  >D��B@  A   >�=q?�K�?�
>��y?Z��D�  ��t>p��D�@ >C�=�oB\)G,mBd(�@�  =�E�G!n�G%�>\(�>�33@\��@�  >�(�>   E��ƶ�oŖXZ?NV   >�bN   A  B�  >�bN=�PE�A��|G@�  >\(�B��qC  D�  ?�/F�>�Ew{�F�z�Dk�ZƲT�E�:�F$�jū�5� D.C�4ř�TƁ'�D�}kF��E����d�A�'uF�zC����v�_E8�ƴ���m����E��-ƃ��Ź��F�D
�NF�2�D��M�u�FŃkF�
��
��F�O��Ÿ���F�Aj�L       split_indices[$l#L       a      	                          
               	            
                                                 
                           
                                                                                                                                                                                                                 L       
split_type[$U#L       a                                                                                            L       sum_hessian[$d#L       aF�` F`P E1� B�  F_ B�  E+  BH  A�  @�  F^� B�  A  E"� C  A0  B  A�  A  @�  @   Cɀ FX� BH  B<  @@  @�  E
 Cƀ C  @@  @�  @�  A�  A  A0  A   A   ?�  @@  ?�  Cg  C,  A   FX� B  A�  AP  B  ?�  @   D�  D�  C�  A0  @�  B�  @@  @@  Ap  Ap  @�  @�  A   @@  @�  @@  @   @�  C9  B8  B  C  @�  ?�  E�  E�� B   ?�  A`  @@  @�  A   @�  A�  D�@ @�  C̀ D!@ C�� A�  A   ?�  @   @@  B<  B�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       97L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       EA��@��YG8�C�]���	�GL~��� C���()���E�C�zF��pE��4�^��E4hgC�*�F��
���LL1�֋]E���nb�G�ƢD�d���1	yF���~\�ů��F��c,��i]F��*�i���@�HeLG�'�F��B��EE��{F���tr�F)���V�yF#���:������kE�w��c�2E]m�Ŧ�<F���ŉ�Í	
F�6D��Ɔ�_�@e�F0M�D��f�1iDE��Ŏ�QD��ƵF��wy�F`�9L       
categories[$l#L                    
          L       categories_nodes[$l#L                L       categories_segments[$L#L                             L       categories_sizes[$L#L                            L       default_left[$U#L       E                                                                L       idiHL       left_children[$l#L       E               	                  ����������������                  !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A����   C������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       EP��P�qOƉ P�(FQ(��O5NP��KQ%�ZPϰ�Q�)�                PQ��Q7\�P��Q��QM)KQb��Q��Q:��Q�`CQ��QS�OQ�zP���P�UzQ4|mQ�3+Q�eyQ�pIQC��Q+PQ_|    P�j,                                                                                                                        L       parents[$l#L       E���                                                           	   	   
   
                                                                                                                 !   !   "   "   #   #   $   $   &   &L       right_children[$l#L       E               
                  ����������������                   "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B����   D������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       EA�     A�  B�     A�  B�33B�  =\@j=qA33F��pE��4�^��E4hgB�  >���B�  ?�@S�
>\)@�\)A��B���=�P=�
=@I�B\��   >hsBY33@N�R@   =aG�@�  A   BP  G�'�BHB��EE��{F���tr�F)���V�yF#���:������kE�w��c�2E]m�Ŧ�<F���ŉ�Í	
F�6D��Ɔ�_�@e�F0M�D��f�1iDE��Ŏ�QD��ƵF��wy�F`�9L       split_indices[$l#L       E                                                        
                                                                                                                                                                                           L       
split_type[$U#L       E                                                                  L       sum_hessian[$d#L       EF�` F�P A   Fg� E  @�  @@  Fc� Cp  D�@ C�  @@  @   @   ?�  F_t C�� B\  C9  D�@ C�  C�  A   FZ  C�� B�  CT  A�  A�  C!  A�  D�  B�  B�  Cy  C�  B   ?�  A  FWP C4  A�  C�  A�  B   C	  B�  A�  A   A�  A   BL  B�  A@  A@  D�@ A`  A�  B8  AP  B�  CZ  A�  B$  Cu  AP  A�  @   @�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       69L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       [A�3��uB��.�T�rGQ��D�x'÷��ŵ�!ǝ�}��� GR�E*��V"F����UFX����:���(�ĭG ��\F��G#��E�E?��+ǞG���E��6��l-D�E�s�G�Q��ē�Ve`��c�<��E����o��F5�E-�Ƌ26G����^��E�"QGbpwD�&���pDŏ<�G3�xFt#�E a�F���č��Ɯ�E�	��y�`F~��CZ�G��FA�qF`�4Ŷ����,z���`�r�F��G\�cE�ZhD�����F��D��U�.gF�X+�+�XE
r���ƅ�rE�A��jF�C�� E��tD�H7�@Q����MCOýD,�_�d^=EWė���&��0CE��L       
categories[$l#L       .            	   
                                               	   
                                     	   
                           	   
      L       categories_nodes[$l#L                            5L       categories_segments[$L#L                                    	       
              %L       categories_sizes[$L#L                                                        	L       default_left[$U#L       [                                                                            L       idiIL       left_children[$l#L       [               	               ����                     !   #����   %   '   )   +   -   /   1   3   5   7   9   ;   =������������������������   ?   A   C   E   G   I   K   M����   O   Q����   S   U   W   Y������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       [Pl�QP]+Q`��Q~��P�ќPc�QF��P���O���    Q!�vQ0�Q\�LP[4"Q)�P��Py�Nr��    L"�QZI�Q88P�M�Qe9$Q8��P��Q>%CQ0�P��OY Pd8�P���                        P�AQѩ�Q��Q�V�PR� P��Qb?Q\v    N}l`P�H[    Q8]Q�x�Qj�GQL\J                                                                                                                                                L       parents[$l#L       [���                                                           	   	                                                                                                                                   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   0   0   1   1   3   3   4   4   5   5   6   6L       right_children[$l#L       [               
               ����                      "   $����   &   (   *   ,   .   0   2   4   6   8   :   <   >������������������������   @   B   D   F   H   J   L   N����   P   R����   T   V   X   Z������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       [<�h@�  >"��B���?L1   =e`B?�Z>�z�@�  GR�@   D�� =�l�>��yD�@ D�� D��    ��\      ?���>���=��   ?}�->��/>�=q?��R   =�9X>��#��c�<��E����o��F5�E-�>�(�>���>;dZ?���B(��@   =��-?/�G3�xD�  ?%`BF���>fffBZ     > ĜF~��CZ�G��FA�qF`�4Ŷ����,z���`�r�F��G\�cE�ZhD�����F��D��U�.gF�X+�+�XE
r���ƅ�rE�A��jF�C�� E��tD�H7�@Q����MCOýD,�_�d^=EWė���&��0CE��L       split_indices[$l#L       [               
       	                         	                                          	   	                                                                                                                                                                                                                                        L       
split_type[$U#L       [                                                                                    L       sum_hessian[$d#L       [F�` B�  F�h B�  A  E� FFD B�  A0  @�  @   EU� Dq  CF  FC, Bl  B4  A   @@  @�  @@  A�  ET@ D� Cހ A   C<  E�8 E�  B\  @�  A�  A�  @�  @@  ?�  @   @   ?�  A   A�  D�� D�� A   C�� B�  C�  @�  @�  C:  @   Eð C  D�� E�� @�  B@  @   @   @@  A�  A  A@  @�  @@  @�  A@  D�@ D_@ B  D�  @@  @�  C)  C�  BL  BH  B�  C|  @@  @@  C0  A   D�  E�� B�  B|  DI  D2@ DT� EhP L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       91L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       }A�YDP��� ��C1޶F	�������D6��Ƴd�FwN7��F��	����+�CZ���E���D��U�#�vFU��G��F�S���ܔĔ�gG�s�Ư�ŔѓF"��ʠPE�W�ü�Ħ.F2�eE�m��:�Gw�3�$.J�%��z�Ť�ZF�ӗG�M�E� 0G�b�FC`�=��F���Gq<��<�G9�Gq�Ƈ��Ǔ؜Ɖ��D`G2��V���|�!��Fg�Ɓ���z� E�O^Dj��JI�G[�nE3�EM���ֆ��Z DǘECIkGC_uŚ�FlF�E|h,�6������(D-ŐêFg�F���E��2F)|�Gj��R�E��`F�G'��F�p�Sm���Zw�F�ڕ��~�F��GE����<�Ù����u:F��mż��F�:^E=����QƔ���l��ĩ��E�H:E�;�F�*�E����'ð��Ɣ��'`�Fkr�C�zE���Ê��ƛ����·��E��=ì�L       
categories[$l#L       3                          	   
                                  	   
                                  	   
                               
            	              L       categories_nodes[$l#L       	                  %   )   .   /L       categories_segments[$L#L       	                                    $       -       0       1       2L       categories_sizes[$L#L       	              
                     	                            L       default_left[$U#L       }                                                                                                        L       idiJL       left_children[$l#L       }               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a����   c   e   g   i   k   m   o   q   s   u   w   y   {��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       }P
p�Q��P�;pQ���Q|܈P��P���Q��Q��rQz�BQɓtQ��P�0�Q�6�P��mQ(+�Q�WQM�aQ���QP5�P޼,Q���Q��P�iSPIܬP�zQ�lQM�Q6lJQQ�P�"Pݪ�Q���Qd
Q�˫Qn7P���P��;Q�jQl��Q�ݮNS NE �P9��Q?^TRֽQ_Nx}�O�2�    P9�P�fJP���Q�Q ��Q�)Q_�Q��^Q�ϖQ,1Q��'P��Q�x�                                                                                                                                                                                                                                                        L       parents[$l#L       }���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <   =   =   >   >L       right_children[$l#L       }               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b����   d   f   h   j   l   n   p   r   t   v   x   z   |��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       }>N�>���=�j>�bN   =y�#>W
=>hr�>D��A�  =�
=BP��>C�D�� =��A33A   >C�B5\)?rn�   >�1@�      =�9X>��#>!��>�hsB�ffB���   D�` >ۥ�>��B�  >>v�   @   ?#�
?�|�   A�B9��@���@ �9      >�t�G9�@��@c�FA   >e`BA�  BI��BVff>)��@�=�/D�` >M��>���Dj��JI�G[�nE3�EM���ֆ��Z DǘECIkGC_uŚ�FlF�E|h,�6������(D-ŐêFg�F���E��2F)|�Gj��R�E��`F�G'��F�p�Sm���Zw�F�ڕ��~�F��GE����<�Ù����u:F��mż��F�:^E=����QƔ���l��ĩ��E�H:E�;�F�*�E����'ð��Ɣ��'`�Fkr�C�zE���Ê��ƛ����·��E��=ì�L       split_indices[$l#L       }                                                      	                              
   	                   	                                                                                                                                                                                                                                                                                                                                                 L       
split_type[$U#L       }                                                                                                                    L       sum_hessian[$d#L       }F�` E� F8 E� D� D=@ Fd E�h C'  C΀ C1  B  D4  C|  Ft E�h D�  B�  B�  Cɀ A   B�  B�  A�  A@  B�  D� B�  C  D+� E�p E�H C�  D�  C׀ A0  B|  B  Bl  B�  C�� @�  @@  @�  B�  B�  B   @@  A�  @�  A   B�  A  C/  CՀ A�  B�  B�  B\  D  B�  E�� D-� D�  Ei @   C�  D�@ C�� B�  C�� A   @@  Bh  @�  A�  A   A�  B  B�  A�  A�  C�  ?�  @�  ?�  @   @   @�  B8  A�  B�  @�  @�  A�  @   ?�  @�  Ap  @@  @�  B�  @@  @   @�  A�  C  C�� B�  A�  A0  B,  B  A�  BX  B  A�  C�  C�  B�  A�  D@� Eè C]  C� L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       125L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       eA�CB�	����jĨ7�C� ��2��-5mE����*1KEi\���Ƨ�E�}��S�K�\3	EO��G�ő�E
�E�3��h}�����D_��F�>N���fŖ�G$�KŜ�ƥ�PE����*��GU�E��'�sw�uʒ�:��F���GMWE�c���#)Ƽ���7������hzE��G=�S�:χƔ*ǒ���I�qF��pG90U���A�(\FEE�E�Dŏ�ů�>F	��F��1E;$ZŒ�[F;vb�.�C�U5�Bk��D��DC�bŻY>Gh.E�ZdFX��żT�EZ������j	dF1���`z�Ƣ0dE��䴕���Ĕ3E�6�ć�
�U̼D�F{F�EZ��� xF%�ś�4��ˀC��N�$�F�h�E�F�$C�q łKE�Y�L       
categories[$l#L                      	                               	   
                     L       categories_nodes[$l#L             	   
            -L       categories_segments[$L#L                                                         L       categories_sizes[$L#L                     	                                   L       default_left[$U#L       e                                                                                        L       idiKL       left_children[$l#L       e               	                        ����            !   #   %   '   )   +   -   /   1   3   5����   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W����   Y   [   ]   _   a��������   c����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       ePLhP��P���P�B�P�W;P��Q{�"P���Pɇ3Q,P��WP�N�P�k    O��~P��P#;�QI�Q1 �Q���P�'�Q2�Q�~P"ϐPp�P���O�$OX��    Pe#�P�؎O���O�,)Q$Q<nQ&�CQ���QjpQ6jP��P���Q	QO��Q*^�QQ�M�`    P��N�* P�kO���O�P        O;!                                                                                                                                                                                        L       parents[$l#L       e���                                                           	   	   
   
                                                                                                                             !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   /   /   0   0   1   1   2   2   3   3   6   6L       right_children[$l#L       e               
                        ����             "   $   &   (   *   ,   .   0   2   4   6����   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X����   Z   \   ^   `   b��������   d����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       e@?+>!��B�(�   >Xb@�p�B�  Ap  ?�bN      @L(�   �S�K@�z�?�Ĝ=�S�?j=q>��T?\(�   >�33>��yB�     @�  @�  @Qhsƥ�PB�  ?�XBz=q>@�?�  B�  AP  >��A  A�  ? �D�@ D� ?%�=�wD�`    �:χ@�ffD�  @��H@ۅD�� ���A�(\F@@  E�Dŏ�ů�>F	��F��1E;$ZŒ�[F;vb�.�C�U5�Bk��D��DC�bŻY>Gh.E�ZdFX��żT�EZ������j	dF1���`z�Ƣ0dE��䴕���Ĕ3E�6�ć�
�U̼D�F{F�EZ��� xF%�ś�4��ˀC��N�$�F�h�E�F�$C�q łKE�Y�L       split_indices[$l#L       e      	          	                                   
   	                   	               
                                              
                                                                                                                                                                                                                               L       
split_type[$U#L       e                                                                                              L       sum_hessian[$d#L       eF�` F�P C  EY FT\ B�  A�  D&@ E/� E� F2� B  B�  @   A`  D!  A�  D�� DF@ D�` D� E� E�� @�  A�  B�  A�  AP  ?�  D
� B�  AP  A   D�� C�� D-  B�  B�  D�� D	� B<  Ee DT� E	� E�� @�  ?�  A�  @�  B\  AP  A�  ?�  @   A0  D� B   B�  A`  A   @@  @�  @@  D� D�  C�� Bp  D� B�  @�  B�  B�  A�  D@ DP� D  Ap  B  A  D� EC  CK  D!� C  E � E!� E� @�  ?�  A�  @   ?�  @�  B  A�  @   A0  AP  @@  @�  @�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       101L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       sA��C[���$��BK�E��ąt	ƊC�B��e�~A�EV��GѧFŎMF0�Ĵ�j�HBFj"�Ǧ�OE��F<��ł6 H;��m����Ʊ�EG�E-T���0UG��P�pN�F���èZ(D�����\G$��˨��	�=G�����l�6�Fژ�B�]�]�FzR�Gtb�Ea�����*Y�E
���(��G61�F���G��F��s��l�:J�G�pF�ŴD�PG�ǞSMŮ�G�3@C!�}ċ��\oBD��6�1���Fj��/�Ğ������ao��~��GϜ�&��E��ƒ �,T�ƫ>�F�6�E��`�D��F;����MŢl�E�x{C�k(F��E��ƒ��Ge�E�K3���[Fp��G"�vE�Q	Ebv�F���*��E[�e�Y�D�u_Gd0}�3��E 'Ft'��6�� 2+E�� ��l�G��E, 4L       
categories[$l#L                                  	                                                L       categories_nodes[$l#L          
         "   #   %   &   *   2   <   =L       categories_segments[$L#L                                                  	       
                            L       categories_sizes[$L#L                                                                                    L       default_left[$U#L       s                                                                                                    L       idiLL       left_children[$l#L       s               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U����������������   W   Y   [   ]   _   a   c   e   g   i��������   k   m   o   q����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       sP�1PWHP�� Ps(Q��Q/�Q.YP�w�Q��~P�A�QſxP�q�QM�~P��Q���P*�rQ��fQU�Q��(Q��QR�O.* N�h�P��UQ�X�QOA�Q[�^P��/O���Q��pP���Q_Q9��Q�3\Qh�P�P�4�Qv��QWo�QB,cQ�&`QDI�QOn�                QWx3P���Q�k�Q�Q�QT��Q@�ZP��Q�3<P�R�Qd�H        O5��P���O��<P��                                                                                                                                                                                                                L       parents[$l#L       s���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   ;   ;   <   <   =   =   >   >L       right_children[$l#L       s               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V����������������   X   Z   \   ^   `   b   d   f   h   j��������   l   n   p   r����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       sA�B�  B��B�  A\)B�ff@�  B�  >��>�hs   B�  @   B   @33@ ��>$�A�  >Z�?��@�        >�S�@�  A@  >E��@@  B  >vȴ@�  @��@��>O�      @�        @u�@�  >��   FzR�Gtb�Ea����A   B}��>]/   >�XA�@�  >�^5D�� B�  F�ŴD�P>49X      B�ffC!�}ċ��\oBD��6�1���Fj��/�Ğ������ao��~��GϜ�&��E��ƒ �,T�ƫ>�F�6�E��`�D��F;����MŢl�E�x{C�k(F��E��ƒ��Ge�E�K3���[Fp��G"�vE�Q	Ebv�F���*��E[�e�Y�D�u_Gd0}�3��E 'Ft'��6�� 2+E�� ��l�G��E, 4L       split_indices[$l#L       s                           
                                                                
                                                                                   	                 
                                                                                                                                                                                                                         L       
split_type[$U#L       s                                                                                                        L       sum_hessian[$d#L       sF�` Fy� D�` Fr4 C�  D�@ B�  FqD Bp  C� A  DV@ Cq  B�  BD  Fp B�  AP  B<  C`  C  @�  @�  DA  B�  Bd  C8  Bt  @@  B  AP  FJ E  A�  Bd  @�  @�  AP  B  B�  C  Cm  A�  ?�  @�  ?�  @@  C�  C�  B�  A�  B$  A�  B`  C   Bh  @@  @   ?�  @�  A�  A   @@  F \ E&� D�� D�  @�  A�  B@  A  @�  ?�  @@  @@  @�  @�  A�  A�  B�  A0  BT  B�  A�  CY  @�  A`  Ch  B8  C� @�  Ap  BL  @   A�  A�  A�  A   A   B  A�  B\  B�  A�  B  ?�  @   @@  @@  AP  A�  @�  @�  @   ?�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       115L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       mA�9(C���� wơ+qC��E���ŀkoĜu	�(�O�DحD�.�D�g�F�Mŝ��F��PF1�����[w�F�K�G\2b�U�D��G �F�6�E�).GfN{E��|Ņ^�@�G��DFy��dw GA��D��@�8j�ǝ�;Ƈ#|E��'D�ŋ�G�$Ơx��&mB"�E��hE�BƦ}�Fz�Ƙ2�G ��,� FȦh�x�_E�l ��ǔ6��H��F,HG
*G6�*B�6�E���d���XgF�"�Ehm����q�!�k�MD����8E����%��E��]�7�G.SF�'�1:�Ɩc`F#�Å�.C�X����iE��nC�~�ź��E�?����Fچ|E���Ď���H���jsEF�����Ǝe#E[)��~2�E��Ɗ\���j��"�$� >�F�	�p�F��OƓ%���S�F� @L       
categories[$l#L       ,                                              	   
                                  
                             	                  
      L       categories_nodes[$l#L       
                         !   )   ,L       categories_segments[$L#L       
                                                  !       "       $       %L       categories_sizes[$L#L       
                                                                      L       default_left[$U#L       m                                                                                                L       idiML       left_children[$l#L       m               	                                    !   #   %   '   )   +����   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G��������   I   K   M   O   Q   S   U   W   Y   [   ]��������   _   a   c   e   g��������   i   k������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       mP#��P���P��3P���P���QpQ0��P%B�P�:�P���Q��P���P���Q_*�QP6_LO�-�P�w�M�
�P��eP�|>Q)�    P�4�P�ڞPj�pP���Q6�Q�I�  P���O|KO���M��'M~��O� O�T�        O^^O�� P��Q2��P�'Q��VP�=P��6P���P/�~P,#x        P�8�Q��?Qp:P�$P���        P���P-d�                                                                                                                                                                                                L       parents[$l#L       m���                                                           	   	   
   
                                                                                                                                   !   !   "   "   #   #   $   $   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   4   4   5   5   6   6   7   7   8   8   ;   ;   <   <L       right_children[$l#L       m               
                                     "   $   &   (   *   ,����   .   0   2   4   6   8   :   <   >   @   B   D   F   H��������   J   L   N   P   R   T   V   X   Z   \   ^��������   `   b   d   f   h��������   j   l������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       m   D�� B0     A@  B(��?c�
>x��>�?�R?�Q�>S��   ?WK�   @33   @�  D� >��D?��By33G �F>z�   @�     >�n�B��B@��?�9XD�  @�     B��A�  BY33E��'D�@�  >�{   ?��R>���   =��
>Ƨ�>t�j>��7?mV�,� FȦh>p��=�\)>�"�@@  B�  F,HG
*?O\)@�  E���d���XgF�"�Ehm����q�!�k�MD����8E����%��E��]�7�G.SF�'�1:�Ɩc`F#�Å�.C�X����iE��nC�~�ź��E�?����Fچ|E���Ď���H���jsEF�����Ǝe#E[)��~2�E��Ɗ\���j��"�$� >�F�	�p�F��OƓ%���S�F� @L       split_indices[$l#L       m                         	         	                             	                          
                                          	                    	      	   
           
      
                                                                                                                                                                                                                    L       
split_type[$U#L       m                                                                                                   L       sum_hessian[$d#L       mF�` Fg� E  BL  Ff� D@ Dޠ A�  A�  EԈ E�P D� BH  Dנ B`  A�  A   A�  @�  @�  E�P E�8 @@  C  C�  A�  A�  D�  A�  @�  BP  Ap  @�  @@  @�  A0  A   @   @   @@  @�  B�  E�P E�� E� B�  B�  C�� B4  A�  ?�  @@  A�  C�� D�` A�  A0  ?�  @@  A�  B  @@  A@  ?�  @�  ?�  @   @�  ?�  ?�  A   @@  @�  @   ?�  @   @   BP  A@  B@  E�� E�( D-  D� D�` A�  BT  B�  ?�  Cl  B�  B  A  A�  ?�  @�  A�  C,  C�� A�  D�� A  A  @@  A   A�  ?�  B  @   L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       109L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       A�EXC�9���E��3�F)�E:#���!C�Ÿ=F� ��'�İ��F]":DU��M��B=9�F+cHFϙ$�6=�F�G3��ƌz�F���E��y�Rg�G$h�E��lF��*ſJ�F�� Ƈ�OC[.*�B��G�?�E�̶�B��G�_�'�������FV��EU
�G��8F�]ƹB�G��%�G��^E���F�,��}��HrsF��&F]OƑ��G[��E4��F�LC�}�Ga7�ƄP��ۗ�E� �@T$�D�_$Ŷ.F)�NG�TFF�3E؈a�TKu���ũ�aF_����8ŋ/�E�,������@�
��}�E/5�E�'��Վ�E��P�s� F��lE���F�!T����B�{�F�;:E�O F3ŴƤ�`FnAF���B�I�E�C)F�bD�C�w����ł@G=n�F�&���IpE����P�IE�Q�FҹwD��]Fv����<D�F�:�:{�Ȼ�F	�GG&�<�����Eş��Ɛ-��ס�F8(\L       
categories[$l#L       ?                      	                	                                    	   
                                 	   
                                  	   
                     
                       L       categories_nodes[$l#L                
                  &   -   =   >L       categories_segments[$L#L                                    	                     '       3       ;       <       =       >L       categories_sizes[$L#L                                                                                           L       default_left[$U#L                                                                                                                 L       idiNL       left_children[$l#L                      	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c   e   g   i   k   m   o   q   s   u   w   y   {   }����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       P�LQ'�Q/YPd8�Q��Q8�QK�PH�lQ�uBQ���Qh,Qm(6Q~�7Q��gQ���P��CP��DQA�Q�Q[��Q��:Q	�P��P���P愠Q��!Q*ʋQ�~jP�EzQ�8Q��P:��Qp�VO��XP�P�Q-fQ/GP
�Q��&Q��HQ��Q��Q#�P���P�Q�P���O8�P��POC�P�EVQP��Q��QG�Qk��Q�EQϚ�Q7��Q�Q�,�Q�Q�(�Qcg\                                                                                                                                                                                                                                                                L       parents[$l#L       ���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <   =   =   >   >L       right_children[$l#L                      
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d   f   h   j   l   n   p   r   t   v   x   z   |   ~����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       D�� D�` @@  D�@    B0     A�  >   B�\)         ?"�>oA0     ?���B�  ?��?�$�>/�@�  >�Q�A�  =���@E�   @�\   @�D�  >�t�A0  >���@�  @IG�B�\   @�  @���>ٙ�?
��D�� ?y��   >��@   ?�\)>�1B�>   >���?��?�(�>�~�D�� A   >L��B��qBL(�      @T$�D�_$Ŷ.F)�NG�TFF�3E؈a�TKu���ũ�aF_����8ŋ/�E�,������@�
��}�E/5�E�'��Վ�E��P�s� F��lE���F�!T����B�{�F�;:E�O F3ŴƤ�`FnAF���B�I�E�C)F�bD�C�w����ł@G=n�F�&���IpE����P�IE�Q�FҹwD��]Fv����<D�F�:�:{�Ȼ�F	�GG&�<�����Eş��Ɛ-��ס�F8(\L       split_indices[$l#L                                                    
                                                                  
                                           
                  
                                                                                                                                                                                                                                                                                         L       
split_type[$U#L                                                                                                                          L       sum_hessian[$d#L       F�` Fk� E0 Fb� D@ D{@ D�� F[� C�  C̀ C*  D4� C�� D� D� FZ B�  B�  C�� C�  B�  C
  B   C�  C�  B�  CY  C  C�  B�  D � FW$ C<  @�  B�  @�  Bh  C�� @   A�  C�  A�  BL  Ap  B�  A�  @�  @�  C�  A�  C  A@  BX  C   Bd  B8  B�  A�  C�  B   B   C�  C)  FMd D  C%  A�  ?�  @�  B\  BL  @   @�  BH  A   C�  BL  ?�  ?�  A   A�  C5  B�  A�  A   B   A�  A  @�  B�  A�  @�  A�  @   @�  @   @   C�  C  @�  A@  B�  C)  @   A   B,  A0  A`  C  B  A�  A�  A�  A�  Bh  A�  @�  B  C�  A�  @�  @�  A�  C�� B�  C  B  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       127L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       qA�\��)��D5?�D�	���;���;EFnUEa��O�Dy�	��T1��ȿǍ/E���Ŵ5�E>�#F�	��e��G�'8EJ(1�#�N�c�nļ�4�gV��l�������E��A�9;���qƜa�EZGB�J�NE�hHQ,FG�Vř��FS� G)ԧń�E�*=Ɣ�DE�����RT�O���ߟ4E�3+F�lc�K5�ŀHmD��fFנSE�}ŵ��F� œ��Fє&���F�
�EIȰC��F�'������FGVPG�_X�W^�D���F�(��8��Q��E�M�E
VI�L+7EyN�ď�#ļE��,P�F3li�!x�E����#�E�w�2ȈĈ����E�L���k�F��Ŧ��0���9W�DR�M�:�wC&ҼF=4FKt�đ�[D�9�E��bYD��"�:qE��x�D�RD��xFO1�E(W��I|��7��F�\��8��L       
categories[$l#L                         
                      
            	                  L       categories_nodes[$l#L                                %L       categories_segments[$L#L                             	                                   L       categories_sizes[$L#L                                                               L       default_left[$U#L       q                                                                                              L       idiOL       left_children[$l#L       q               	                                    !   #   %   '   )   +   -   /   1��������   3   5   7   9   ;   =   ?   A   C   E   G����   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c   e   g   i   k   m   o������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       qO�s�Pҵ�Q:P�Q(��Q���P�YdQ@��QOQ!b�Qw��Q�p0P�<O(ǠQ/��P�8�Qn)�RVP�LP��Qe|TQZ��Q�vQOz�Q>�NP��        Q��Q���Q ��P��Q9M�R#�Q��[QɋP���P��\NH�    QSo�Q�ǿQ��Q� Q�/�Q&h�QW$�Q���Qv}P�n�QN�Q3ޜQ8*�Q#1�QJ�^Q^�DP��P)��Pǯ�P�s�                                                                                                                                                                                                                        L       parents[$l#L       q���                                                           	   	   
   
                                                                                                                             !   !   "   "   #   #   $   $   %   %   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   :   :L       right_children[$l#L       q               
                                     "   $   &   (   *   ,   .   0   2��������   4   6   8   :   <   >   @   B   D   F   H����   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d   f   h   j   l   n   p������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       q   @@  @@        C     B���AP  D�� B�ff   B�B���   B���@�  =���>	7L? Ĝ?Z>H�9>���>k�?\j�������D�  B�  ?��H   @	��@   >,1A@  >�Z>Ƨ�   G)ԧ=Ƨ�>�-?���>� �=�hs>t�j>��\>�!D�  >�o>333BfffA�  @�  @J>���B���@�  ?w��@�  EIȰC��F�'������FGVPG�_X�W^�D���F�(��8��Q��E�M�E
VI�L+7EyN�ď�#ļE��,P�F3li�!x�E����#�E�w�2ȈĈ����E�L���k�F��Ŧ��0���9W�DR�M�:�wC&ҼF=4FKt�đ�[D�9�E��bYD��"�:qE��x�D�RD��xFO1�E(W��I|��7��F�\��8��L       split_indices[$l#L       q                                                                           
                                                                               
                  
         
                                                                                                                                                                                                                           L       
split_type[$U#L       q                                                                                                         L       sum_hessian[$d#L       qF�` FX Fh E�� E� E�� E�@ E)  D�` E!� D�  E�h @�  Ee� D  E%` Bh  D�� @�  EP CҀ DJ@ D�  C� Er� @   @@  E� D�  Cހ B�  E$  A�  BT  @�  B�  D�  @@  @   D7  D�  C�  C  C C�  D$� C�  Bx  CҀ D�  E B�  E� DP� D� C�  B  B�  A�  D-  D�� @�  A`  A�  A�  @�  ?�  B�  A0  D  D4@ @   ?�  C�� C� Dc� D� C  B�  B0  B�  B0  C�� B�  C�  D� B�  C6  CX  B,  A�  B8  C�� D  D9@ E� B�  B�  B  DР C�  D� C�� C"  C�  C�  C  A�  A�  BH  B@  @�  AP  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       113L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       UA�~�B����%�aC�^����#�`���)RC�� ө�lo5�Х�F_�^ܰEb�Æ�Z����8BmC��{�@���a�G>��FaTEt�ƥ�&F,�B��:F��C��ŉf��#(�`YfF�,��;[hĎ��F_mƏ=�ƨ��?W4F�pGj��F�Թ�_l�F.�D���#���w�/ F1�MFTF��a�~�	n�E�aEܞB�����o�/��ż�F�q��&/�/|�E���F�nE��&��I�D�gj��ͭFj��D{�D���:4�%���R��D*�F�(��ɫF0��Cw\ūo'��^�E��}Eu�M�)�����uE�@�ų2�C��4L       
categories[$l#L                       
                          L       categories_nodes[$l#L                      *L       categories_segments[$L#L                                           L       categories_sizes[$L#L                                          L       default_left[$U#L       U                                                                           L       idiPL       left_children[$l#L       U               	����                                    !   #   %   '����   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C����   E   G����   I   K   M   O   Q   S������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       UO�j�O粙O�_�P�m�P�Y    O�(P��NP�N�P���Q|N��6O�XQ��qP� �P�VdQ]�Q�dP�hQb@QK|L    O�!O�2O�rdQz Q�`fQ��Q��P�EPYN�P�)�Q(v�Q��Qs0$O~��    Q4�#Q��    P,��M��~MՑ�O��O�0tNF�                                                                                                                                                            L       parents[$l#L       U���                                                     	   	   
   
                                                                                                                                   !   !   "   "   #   #   %   %   &   &   (   (   )   )   *   *   +   +   ,   ,   -   -L       right_children[$l#L       U               
����                                     "   $   &   (����   *   ,   .   0   2   4   6   8   :   <   >   @   B   D����   F   H����   J   L   N   P   R   T������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       U@��;   =�x�B�     �`�   @=p�=�h@�Q�A33>Ǯ   B�  B�  ?!G�>@�@���A   >�ȴA��FaT@   @@  B���<�t�>fffD�` @XQ�Btp�@�  >�ƨB�R@@  @�\)?G�ƨ�>�bNA�  Gj��@   @@     D�@ D�` @�  F1�MFTF��a�~�	n�E�aEܞB�����o�/��ż�F�q��&/�/|�E���F�nE��&��I�D�gj��ͭFj��D{�D���:4�%���R��D*�F�(��ɫF0��Cw\ūo'��^�E��}Eu�M�)�����uE�@�ų2�C��4L       split_indices[$l#L       U   
                                                                                                 	                                                                                                                                                                                                        L       
split_type[$U#L       U                                                                                L       sum_hessian[$d#L       UF�` F�� B�  Ff� E @�  B�  Fb� Cp  D� D  A�  B<  EP F# B   CH  D�� Ap  D@ A0  @@  Ap  B  A0  EC� Dn  F
p D�  A�  A�  B,  C  D�  C&  A   @�  C�  B�  ?�  A   @�  A0  A�  AP  @�  @�  A�  EB� C~  D.� B�  F	< B�  D�@ A�  @�  @�  Ap  B  A   B8  B�  D/� Dh@ B  C   @�  @�  C�  B   B�  AP  @@  @�  ?�  @@  @   A  @   A�  @�  @�  @�  @@  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       85L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       /A�B�@�2�G�{F����+���w��G^� G_��3�7�!��C������DF(�F�o�E�ޚ��f�GB�_E�&���E���A�jF���E�v'�7ʡF����	l;FF/�G�DY ��x~6CyiĬ�F�wFMy��&��P��ś��E�HE�q��FU��ś��E�����q_����W�E��?Bq�oL       
categories[$l#L                                      	   
                L       categories_nodes[$l#L                   L       categories_segments[$L#L                                    L       categories_sizes[$L#L                                   L       default_left[$U#L       /                                          L       idiQL       left_children[$l#L       /               	         ����      ��������������������               ��������      !   #   %   '   )   +   -����������������������������������������������������������������L       loss_changes[$d#L       /O��O��]PX�P!�O�sNo�N:`O�ת    P�
4PG��                    N`��Q>}P�Q,�KPQ�        P�\rQe�Pڰ(Q4pP��DPԠyQ:�P�S                                                                L       parents[$l#L       /���                                                     	   	   
   
                                                                              L       right_children[$l#L       /               
         ����      ��������������������               ��������       "   $   &   (   *   ,   .����������������������������������������������������������������L       split_conditions[$d#L       /CJ  D�  D�@    ?=p�B�33   >����3�7>^5?>o����DF(�F�o�E�ޚ��f�>�C�>:^5A0     =49XF���E�v'B���>߾w>x��   B�  =�9X=��?E�Ĭ�F�wFMy��&��P��ś��E�HE�q��FU��ś��E�����q_����W�E��?Bq�oL       split_indices[$l#L       /                                                                                        	            	                                                                   L       
split_type[$U#L       /                                           L       sum_hessian[$d#L       /F�` F�T @�  A  F�B @   @�  A   ?�  Dz  F|� ?�  ?�  @@  ?�  ?�  @�  C�  D0  C�  Fx� @�  @   Ce  B�  D@ B�  BH  C`  DO  Fk� CK  A�  B`  A0  C�  C�� B�  @�  B$  A  B|  C!  B�  D0@ A�  Fk< L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       47L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       AkU�D��TÖ�bE��UĠ�IƇW���ED��'F\���F��0F�?���N��n�DE����N^��m��F�1J�}��E�֭Gg�_Cr�G3�sDct��>=���(vC���=��E�9XśL��?��E�18D�ex����C�{�<N\F>o�GA���;��*\KD�k�F�fF��Hq�G��N���VG}^�F�ðƬ�F�2gǥA���"F�FG�3s�D֥��A�;����EH��Ų�oE�C���ӎ����£�����E�Z�D2�<�_4F!o�����(E���j�ưpE�	{E��ų��Fr#F�3���{F�D��(ŪO�Fw��CDw'F�L�2�FUw��tWD|8gGX2`GFD�T�NE`����ݎE��F���F6��ś��E�Z�`WE�p.�ȁ��Ak�"�!�@�FLP�F�@D�mƶ�^ŦD����ԃ}�N�Ɠ��V��D����YگE��F����n~F�D�NV�/E~F�Ý� ܲE38�L       
categories[$l#L       O                         	   
                                  
                            	               
                                            	   
                                            	   
                               	   
            L       categories_nodes[$l#L          
         %   (   -   .   0   5   6   7   <L       categories_segments[$L#L                                                  %       &       '       (       5       6       AL       categories_sizes[$L#L                                                                                           L       default_left[$U#L                                                                                                             L       idiRL       left_children[$l#L                      	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c   e   g   i   k   m   o   q   s   u   w   y   {   }����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       O���Q��Q��Q1ޜP��QK�XP;�FQG��Q���P��QI�.P_bJQ$��P���QC_7P�t�Q�Q��Q��Q�.P�,`Q=��P�0�O��|O��Q�QO��Q��Q�b�Q.Qw��Q*��QCQ&�)Qsb�P#@�Q/Y?Q�#QLrP��CQwl�P�K(Q�zP�ǈP�-�P��PV��M	C�O�%N��O��Q4a
Q�6Q��P�)�Q228Q:��Q���Q��P�c�Q�(�Q�s.Qn"                                                                                                                                                                                                                                                                L       parents[$l#L       ���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <   =   =   >   >L       right_children[$l#L                      
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d   f   h   j   l   n   p   r   t   v   x   z   |   ~����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       >�>8Q�>�9X>�>�`B=��#@���>   =�x�>�      D�@ @��@>�+<D��B  Bh  B�k�>(��B��{?�/>Kƨ@�  >�o   @�  @�  @bND�  @K�
>��=�jA�  >��T>C�>1&�   >��A     >Y�?��BZ  B��      @      B  >���>��H@�           CW
@�  D�� ='�   B��{D�� £�����E�Z�D2�<�_4F!o�����(E���j�ưpE�	{E��ų��Fr#F�3���{F�D��(ŪO�Fw��CDw'F�L�2�FUw��tWD|8gGX2`GFD�T�NE`����ݎE��F���F6��ś��E�Z�`WE�p.�ȁ��Ak�"�!�@�FLP�F�@D�mƶ�^ŦD����ԃ}�N�Ɠ��V��D����YگE��F����n~F�D�NV�/E~F�Ý� ܲE38�L       split_indices[$l#L                         	         	                                                                                                       
                                                                                                                                                                                                                                                                                                                                   L       
split_type[$U#L                                                                                                                          L       sum_hessian[$d#L       F�` E^  FU@ D�@ E	` C  FS0 Di@ CҀ E� B�  A�  B�  F,� E D7� CG  B�  C�  DƠ D  A�  BP  A@  A�  BL  BP  E�� E3� DԠ D?  A   D5  B�  B�  BD  A�  C�� B�  D�� D� C� Bt  A�  @�  @�  B@  @�  @�  @�  A   A�  B  A�  A�  E�� E� D�@ D�  C�  D�� B�  D*  @�  @@  C  D@ B�  A�  B�  @�  A�  A�  A�  @�  Cv  A�  B<  A�  D~� B  C   C�� A   C� A�  B  A`  @@  ?�  @@  @   @   A�  A�  ?�  @�  @�  @   ?�  @�  @�  @@  A@  @�  A�  @�  @@  A�  A  A@  D�� E�H E� AP  D�� C�� Cy  Dz  @@  C�� C
  D�` B�  @@  C� CW  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       127L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       {A��]�X|Cd&�Ş��E�e�E�B��F��ƶ�hE=�jG��FvFƶz3Ũ�C�SFC��ƖI#�8] �<�4�Q�F�0�G�%AE�:��(0@F��������BG:,(���F��kB�%�E����޳�s%x���ƍ*gG�p���\� �|E� ���[jG9�����Fx�`H�AGN�0�v�D��P�FgVG]�jC � F4%Ǐ���ޭEB���6u7G��s�A��Gx���G/��oy?C+��D�XF�����hćg�D4)�ϕ�s6y�^�|G	z�egų�M��)�M�E�d�FZ��B��C��lF��E��?F���űKF0C�E��Z���E��G8�4F��E�;�Fk���Y'��[n�f�}��:�F&@QG
 &F,܇ıU�G(��J�KF�������D�� ƞs��]%vF�8�q��E��YF��MŖ��E�O�F���g�E�E�?rE01F���E��*�4�D�ؘ�B�|�L       
categories[$l#L                               	   
                              
                                      L       categories_nodes[$l#L       	               +   ,   .   /   ;L       categories_segments[$L#L       	                                                                L       categories_sizes[$L#L       	                     	       
                                   L       default_left[$U#L       {                                                                                                           L       idiSL       left_children[$l#L       {               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C����   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c   e   g   i����   k   m   o   q   s   u   w   y������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       {P u4Qv�Pjk�Q\<NQ��QyAEPZ��Q�!Q!\�P�l�Q4��Q���Q�E�Q�O7Q'��Q�Q$�lQb�cQ��Q:G�Q�nPӡ�P��jQ�lQŒqQM�KP�2�P۹�Q��Q�iDPk+�Q/a�QjQ%�    P��BP�&~O��`P��Q"1\P��&QJ`P=N NU�tP�$�ME�P�c�P���P7))Q��QiP�2�O��HOE@    PI��P�1 Q8!Qj`Q���Q��Q>��P*.                                                                                                                                                                                                                                                L       parents[$l#L       {���                                                           	   	   
   
                                                                                                                                         !   !   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   7   7   8   8   9   9   :   :   ;   ;   <   <   =   =   >   >L       right_children[$l#L       {               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D����   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d   f   h   j����   l   n   p   r   t   v   x   z������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       {>49X>e`B>G�>�(�B��=@��R>gl�      >��uA�  B@  D�  =�E�>p��Bb�\?   >� �@�  >	7L   @�  >���D�     A0  >B�\>aG�A@  @@  >vȴB`  Bq33=ě����=��B���B*�R?��>{�mB,  Bq33>��      B�        @�  >z�Ap  D�� B�  B�  EB��@   D�@ @�  B     BL(�?��=t�D�XF�����hćg�D4)�ϕ�s6y�^�|G	z�egų�M��)�M�E�d�FZ��B��C��lF��E��?F���űKF0C�E��Z���E��G8�4F��E�;�Fk���Y'��[n�f�}��:�F&@QG
 &F,܇ıU�G(��J�KF�������D�� ƞs��]%vF�8�q��E��YF��MŖ��E�O�F���g�E�E�?rE01F���E��*�4�D�ؘ�B�|�L       split_indices[$l#L       {   
      
            
                     	   
         	      
                       
            
                	                     
                                                                                                                                                                                                                                                                                                                L       
split_type[$U#L       {                                                                                                                  L       sum_hessian[$d#L       {F�` D�` Fv� D�  C�� C�  Fr� Dn@ C  C�� A�  CV  BX  C�  FkL DP@ B�  B�  B<  C`  B\  A@  A   B�  C  B@  @�  A�  C�  C  Fi, C�� C�  B�  @@  B�  @�  A   B  C  B�  B   A�  @@  A  @�  @@  B8  B  B�  Bl  B  A  @�  ?�  @�  A�  C�  B  Bx  B�  B�  Fh( C�  A0  B<  C�� Bd  Bp  A`  B�  @�  @   ?�  @�  B   @�  A�  C  B�  @   A�  @�  A�  @�  @   ?�  @   @�  @�  ?�  ?�  @   A�  A�  A�  Ap  A�  Bd  Bh  ?�  B   @�  A   ?�  @   @@  @@  @@  A   A   C�� B$  A�  A   A�  B   B   B  A�  B  C�� Fc< L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       123L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       {A���C�yvĴd�B��FF�p�E8M�ŚK!�>!�C�M�F�u��7��F4{��TA�&.��f`�ž�]E�b�Eɮ��jc�e�qG�a��oSFU�{E
�>F���DҊZƶ�?ũ ���oF�XB�CB���2F��ER9GƇ�Ed�G��Cg�������g�ƢX�F��1G��}��'c�l;�;+Gv��E�w��;{�G���F�q�ņ�HF��$E�/�#3���_VG���ǀ�ƌ��G���FH~7��Z��n�ĈηŦzuF�d;D X�_/bE���G)�E���E�r�)��E�m�F��<BcZF�,Ĺ2��lŹ�\FO�Ĭ�4F�9O�
����=B��Ƣ1FxŸ�<F�����~��_GED��FYƋ�T�C?3G<�F&���&0�
 D~�&Fz��B�E�޿�y���@C�?Wô�*�>�ƕG�"F�e��S-D�D��39hG.���M�TFA�������LEN�ZƮ'�E��{L       
categories[$l#L       &                                               
                                              	               
          L       categories_nodes[$l#L       
      
                     *   5L       categories_segments[$L#L       
                                                         !       $       %L       categories_sizes[$L#L       
                                                                      L       default_left[$U#L       {                                                                                                          L       idiTL       left_children[$l#L       {               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M��������   O   Q   S   U   W   Y   [   ]   _   a   c   e   g   i   k   m   o   q   s   u   w   y������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       {O�)�Qg��Q%�eP%�Q�3�Q���Q!v8P� P�9�Q3�8P�j$Q�v�Q�]�Q��Qaf�P���Q�o�Qg<�P���OD��Q-�P���Pֆ�Q��FQ���Qs3�Q�ZSQ���Qnr`Q�G�Q{��P�:Q5�%Q6�PTF�Q��Q"!P^��Q���        P�4VP���M2� P�37PW�PDwQ���P�R�Q�R�Q���Q���Q���Pԧ�Q?xpQ��nQ-�Q��QS�QXլQ(�Qf�kQ�,�                                                                                                                                                                                                                                                L       parents[$l#L       {���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   $   $   %   %   &   &   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <   =   =   >   >L       right_children[$l#L       {               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N��������   P   R   T   V   X   Z   \   ^   `   b   d   f   h   j   l   n   p   r   t   v   x   z������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       {B�  B�aH?j=qD��    @�  ?H��@�  D�  >���   @�  ?:^5   >dZ?o@�  B�        A   @@  @?\)>���A`  ?%`B   D�  @      A      >Y�>��@�  Bh  >_;d@�  @�  �g�ƢX�>,1   B�  @)�#>G�@*n�=�Q�>�P>�X>�
=B��=@@     ?E�TD�� B�  ?�z�D�  ?˅B��{D�` ?��ĈηŦzuF�d;D X�_/bE���G)�E���E�r�)��E�m�F��<BcZF�,Ĺ2��lŹ�\FO�Ĭ�4F�9O�
����=B��Ƣ1FxŸ�<F�����~��_GED��FYƋ�T�C?3G<�F&���&0�
 D~�&Fz��B�E�޿�y���@C�?Wô�*�>�ƕG�"F�e��S-D�D��39hG.���M�TFA�������LEN�ZƮ'�E��{L       split_indices[$l#L       {                      
                  
                                   	                                 
                                         
         
               
               
         
                                                                                                                                                                                                                                                L       
split_type[$U#L       {                                                                                                                 L       sum_hessian[$d#L       {F�` F_p E5@ F\l CA  D�� D�� D�  FK� C
  B\  D@ D9  D6� D]@ DG� C�  D.  FA @�  C  A�  A�  C�� C6  D� C  D� C#  B�  DE@ D:� BT  C{  @�  D @ B\  F:d CԀ ?�  @�  B�  A�  @�  A�  A�  @�  C�� A�  A�  C!  C�  C  Bl  B�  D� A   B  C   A   B�  D6� Bh  D@ C]  A0  B(  B�  C	  @�  @   D  BD  B  A�  F:$ A�  C�  A0  A`  B�  @�  A�  ?�  @�  A�  @�  @@  A`  @�  ?�  A�  C�� @@  A�  @�  A�  B�  B  B�  C�  BT  B�  B(  A�  A�  B�  C�  B�  ?�  @�  A   A�  Bx  B�  @�  @@  B  BT  C߀ C�  B  A�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       123L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       aAd0(�Av�C
��F*'��E��6A%���t� Ņ)e�����9����.Fb:���T�E~j�Ɵ�<�g���T&ǃcEv���飏�a>�G��XF�NH�G
WB�0^ō�HGuE��F��)��RF5+Ǥs�G�	C��E�Mƣ����;E�A�GB�D���GG����ƣ�G2��C������,�7�MfCE��G���Y�F�F���%������+��E�]�D�.��o��#F:F���Ɔ�0�,F�MC11kFf?s��d7�7\�Oy7Ƶ��Ev�=�rE?�Fp#0E���;%-�5+�;�E��;F�A�:�D�j�J�n�q��v�SD���AV��BY]Eޡ1���F�bņ���〳E ��E��+�-H�L       
categories[$l#L                             	   
                                            
      L       categories_nodes[$l#L          	                   !   ,   /   2   4L       categories_segments[$L#L                                    	       
                                          L       categories_sizes[$L#L                                                                                    L       default_left[$U#L       a                                                                                   L       idiUL       left_children[$l#L       a               	         ����                  ��������         !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G��������   I   K   M   O   Q   S   U   W   Y   [   ]   _��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       aOƺ�P�$Pf��Ohw�P�/�Q rmPX�N��     P�ǬP�q�Q#�6Q"E8P^�fP��        PqnP}?$Q)�QxQ�P��Q>�RP�X�P@��Qg�Q	�+P��P�dO��BJhn�P�@Q�tP��P���P�f�Q�/P��        Qw�QU�P	LP1�PsNtP�[QRB�Q�YPY�PS[0Q1%3P�U6                                                                                                                                                                                L       parents[$l#L       a���                                                     	   	   
   
                                                                                                                             !   !   "   "   #   #   $   $   %   %   &   &   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4L       right_children[$l#L       a               
         ����                  ��������          "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H��������   J   L   N   P   R   T   V   X   Z   \   ^   `��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       a=��
=�=ě�=��@@  >1'B�  =��Ņ)e   >JB�     B�  =uƟ�<�g�   @"�\   BW��D�  @�  >��wD�@ @CoB�  ?�y>o��?���>t�j         ?WK�@0A�> ĜB<�H?��`GB�D���>ۥ�B���>�   @�  @�     =�j>���   B     F���%������+��E�]�D�.��o��#F:F���Ɔ�0�,F�MC11kFf?s��d7�7\�Oy7Ƶ��Ev�=�rE?�Fp#0E���;%-�5+�;�E��;F�A�:�D�j�J�n�q��v�SD���AV��BY]Eޡ1���F�bņ���〳E ��E��+�-H�L       split_indices[$l#L       a                                                	                             	               	   
                            
           
                                                                                                                                                                                                                   L       
split_type[$U#L       a                                                                                      L       sum_hessian[$d#L       aF�` D%� F�4 A   D#  C�  F}� @�  @@  B   D  B�  CJ  Fu� C�� @�  ?�  A�  A0  C�� C{  B�  @@  C  B4  Fj� D6@ A�  C�  A@  A�  @   A  A�  C�  C  B�  B  B4  @   ?�  B�  B`  B   @�  FQ D̠ D0  A�  A�  A  C/  C�� @�  A   @�  A@  ?�  ?�  @�  @�  A�  @�  C�� ?�  B�  A  B�  BL  A�  A`  B(  @@  B  Bx  B   A�  A�  A�  @�  ?�  F?� D�� D�  C|  C�� Cʀ A�  @�  A0  @�  A   ?�  B�  B�  Cj  B�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       97L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       E@��U��݌F�w�D��#5��~XG9YC@�FJ@��:�F�K�FD�pC���=r��/L�F�#E3f��x4E5�Ŀ�-¾� E���B���FK#K�9u��/y#G9_őM�GQƧ��FG��D��G��Ɗ�E���Ő�\E+�_�_D�D3�����F��E=��Ɯ�D�Nƴ��ų��.�(F��FN�Cƃ�-���q˷D�o�F1�%ƀ�}D��aG���ԅ�D�+��3E�oDQ��k�E��E����D����ԑL       
categories[$l#L       !                	                        	                         	   
                                    L       categories_nodes[$l#L       	      	                  !   %L       categories_segments[$L#L       	                                                                L       categories_sizes[$L#L       	                                                               L       default_left[$U#L       E                                                         L       idiVL       left_children[$l#L       E               	����               ����                     !   #   %��������   '   )   +   -����   /   1   3   5   7   9   ;   =   ?   A   C������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       EO�[�O�'aO��jP���P�3    O�P�h;Qh��QC�JP���    M^�8Qq�QG�8QCC.Qd�:Q�Q~��Q��Q��        P�͓QuR?Q|�oP�v0    P�YhQ��O#DQ�Q��uP�<�Q �QIV�Q/� Q��;Q%�'                                                                                                                        L       parents[$l#L       E���                                                     	   	   
   
                                                                                                                 !   !   "   "   #   #   $   $   %   %   &   &L       right_children[$l#L       E               
����               ����                      "   $   &��������   (   *   ,   .����   0   2   4   6   8   :   <   >   @   B   D������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       EA�  B[z�D�� BX  Ba���~XA�  BU��      @�  F�K�B��BS�HA   @         =L��      ¾� E���D�� =uD�@ >O�;G9_   A   ?ƨD�  >G�   >+>�7L?�|�   >8Q�D3�����F��E=��Ɯ�D�Nƴ��ų��.�(F��FN�Cƃ�-���q˷D�o�F1�%ƀ�}D��aG���ԅ�D�+��3E�oDQ��k�E��E����D����ԑL       split_indices[$l#L       E                                                                                  	                   
                                                                                                                                                 L       
split_type[$U#L       E                                                            L       sum_hessian[$d#L       EF�` F�P A   F E� @   @�  F  C�� D� E�0 @@  @@  FX C2  C-  C  C�� C�  E@ E�� ?�  @   F� Cs  C  B  ?�  C,  B�  A�  C$  B�  @�  C�� D� C�  D�  EL E�� E�0 @�  Cm  A`  B�  A�  A�  C  A�  B�  A�  @�  A�  B�  B$  A�  B�  @@  @   B�  C  C�  D�� C�  C@  C�  D�� D�� E� L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       69L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       A.j�C�2�ģ���xY5D�c}C�8_��0�D�`,�ĞUŗ��D����\eF����w��D��-EIf���M�v:2ƴcF[P����PE��&D�sE�8�$e�F$kG�q_�qW���qF�ƒ�%FVn�D߁�F��r��AŤ�IF�IN�Ei�ǂ\jG4�D�wŵ-��k=Eѯ>�S��D�F��W�xɩFW)	C��E��G&��E��G��eG��F��[�J��nrlƭ]I�S��F�:�ƽߩF��E���=}D۴����	�	�ZF)��ž� �n��ėg����uF� ��Q5F���Ō-�F����@IŚ؜F�؋Ev�ƅ���SG#�*D�M��LCb7UEz�TƳ�>E���(�D�!�FQ;�c\DL���W{OE,?pF����XC����ْV�-"�F�O�E3#��]�+EL *G#�iE���FOV~De�����F�U	�D���<0������Jź���ЊF�ʧD�:�F��E?������MFm+L       
categories[$l#L                 
                              	       L       categories_nodes[$l#L                        !   (   0   6L       categories_segments[$L#L                                                  	              L       categories_sizes[$L#L                                                               L       default_left[$U#L                                                                                                                       L       idiWL       left_children[$l#L                      	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c   e   g   i   k   m   o   q   s   u   w   y   {   }����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       O���PD�!Qr�QK3P�@Q�gQ5��Qz�8QNLQ��Qe�P���Qr:QY��Q/%Q"x.Q�2QZYfQ���Q(� Q Q� .Q��Ql_P��P���P"�8P��XQ
��Q��P��Q�A)Q�QJm�Q.�HR
��Q�3jP�ciR�P��P�edQm�PQ�.0Qs�fP���P� QM��P���Q���P��P��P�?�P%��O�� N&�Q�UOQE��Q�BP�,P���Q;PW��PBLb                                                                                                                                                                                                                                                                L       parents[$l#L       ���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <   =   =   >   >L       right_children[$l#L                      
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d   f   h   j   l   n   p   r   t   v   x   z   |   ~����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L          @   @�z�@�  =�j@���@	��   D�� =��>(��@      D�� ?�/=�`B=�oB�(�B�  >�-B��?wK�Ap�Bo33Bo33D�� ?G�>z�>-VD�� B�=q@ȣ�      >cS�B��B�
==u?�{>G�   B�  =�t�@��R?�;dD�@ =�o?
��   @@  A0  ?	x�>D��D�`    D�@ @#ƨB{��@�p�A�HBP��D�� ?�7LE���=}D۴����	�	�ZF)��ž� �n��ėg����uF� ��Q5F���Ō-�F����@IŚ؜F�؋Ev�ƅ���SG#�*D�M��LCb7UEz�TƳ�>E���(�D�!�FQ;�c\DL���W{OE,?pF����XC����ْV�-"�F�O�E3#��]�+EL *G#�iE���FOV~De�����F�U	�D���<0������Jź���ЊF�ʧD�:�F��E?������MFm+L       split_indices[$l#L                             
                                              	                                                	                      	                                                                                                                                                                                                                                                                                                                      L       
split_type[$U#L                                                                                                                              L       sum_hessian[$d#L       F�` F[� EC` E�P F@ E� D#� Ec D�  DX  E�� E B�  C�  C�  E5  D8@ D�� C+  B�  D>  DЀ E�` D8� D�� B�  A   C>  C$  CZ  B�  C�� EP Bl  D)� D�` B,  C  B   A�  B�  D3� B(  D�  A�  E�  C�  C�  C�  Du  D� A�  B�  @�  @@  B  C  A�  C  C  B�  B�  A   Cf  B�  D�` D�@ A�  B(  C~  C�  D�� AP  A�  A�  @@  C  @�  A�  @�  A�  B�  A   D3  @   A�  A�  DY� DB@ Ap  @�  Ev� E� A�  C�� C�  B�  C}  A�  A�  Do@ D  A�  A@  A   B  B\  @�  ?�  @   ?�  A�  @�  B�  B�  A�  A`  @   C  C  @   B  A�  A   B�  @   @�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       127L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       sAX_�ud�CḡB��$����Et��TS��tׇC�Hr��0pGƐE�$��92U�P�	Du�E�6�&M��LD�����Gb��G;^zF�0LF[��CH��FO;��	��E2����_E�=�ýF��>šuwǁ�PEg�Ƈv���ΘD�h{GFE����J��G
%jEڬIF���F0��<m,F��mƎ��E��5F�J����U�� ��;P�F�]��T��E�5�H�ER5F���C�����2F��D�FŢ��E�������0�;��Fkf��]%�Ƨ6,ķD��RE.��B�Ȅ�+�=F{=1F��WC����'���4ZFc_gŵ*E��e�P��FA}Ņ��F��mE�9�F�rv�η�ED��Ž� �S@yF`�XƐ��]���"�iFܐ�E e�F<��/��EΎ�C0��Flc%ńr,�U%Dv��3��F2'�ŷI��{�ME	��]�G�R�9L       
categories[$l#L       .                           	                                                                      	   
                                       	   
      L       categories_nodes[$l#L                         !   (   *   ,   .   5   6   :L       categories_segments[$L#L                                                                                     #       $       %L       categories_sizes[$L#L                                                                                                  	L       default_left[$U#L       s                                                                                             L       idiXL       left_children[$l#L       s               	                                    !   #   %   '   )����   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O����   Q����   S   U   W   Y   [   ]   _   a����   c   e   g   i   k   m   o   q������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       sO�h�P�cP��	P�r&Q/MAQ!�\P�0mQʢP�ʞQ5�P��Q%�uQJ��Q�rP���P���QN7ZPؼ�P�<�Q(��P�2�    P��Q)��P�yDQ��BQ�B�QK�P�rQu�PP��P��P h	QYPP,�Q P�A�P��P�nQ+Qc�p    O��H    O���QdjQ�|P���Q3��Q���P�R�Q�D    P�s�P���Q��P���Qb�hQ��>QR0mQ�`                                                                                                                                                                                                                        L       parents[$l#L       s���                                                           	   	   
   
                                                                                                                                   !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   *   *   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <L       right_children[$l#L       s               
                                     "   $   &   (   *����   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P����   R����   T   V   X   Z   \   ^   `   b����   d   f   h   j   l   n   p   r������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       s> Ĝ>\)>C��@   A�  A�  >�   >n�@�  @   ?_|�D�     >u   ?j=q   ?�|�>n�D� G;^z=o>�@   >��@�     >hr�B�33B�  ?>5?@      @�E�@#ƨ?R�!>1&�?=�@@     G
%j   F���   ?��   >!��>ٙ�>�bB  A,���;P�      >A�7>��uB�\   A�  >��uF��D�FŢ��E�������0�;��Fkf��]%�Ƨ6,ķD��RE.��B�Ȅ�+�=F{=1F��WC����'���4ZFc_gŵ*E��e�P��FA}Ņ��F��mE�9�F�rv�η�ED��Ž� �S@yF`�XƐ��]���"�iFܐ�E e�F<��/��EΎ�C0��Flc%ńr,�U%Dv��3��F2'�ŷI��{�ME	��]�G�R�9L       split_indices[$l#L       s                     	                
          	      
                                              
               
                                                                              	                                                                                                                                                                                                                        L       
split_type[$U#L       s                                                                                                      L       sum_hessian[$d#L       sF�` E�@ F:� E�p DN� D�� F"� B�  E�� DH� A�  Dl� D� D�� F� B|  BL  D�` EB DF  A   ?�  A�  D@ C̀ C  C�  D� D�` D�` E� A�  B0  B  A�  C  D�  E@0 A�  C0  D  @�  @�  @@  A�  B�  C�  B�  C�  B�  B0  C�  @   B�  C�  B�  Di@ D�@ CA  E�P D  A   A0  A�  A�  A�  Ap  Ap  @@  B�  A0  D@� C�� Cڀ E$� A   A�  @�  C)  C�  CT  @   @�  A@  A   A�  B�  A�  Cƀ @@  B�  C�  Bx  B  B�  A0  B  Cπ @@  B�  B   C�  A�  B�  A�  D  Cƀ D�� B  C  BX  E�( DI@ Bp  D  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       115L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       }A�U�� D1R�6����śF4[�C��ƨ݁�c�ïE�Ɨ��F�15���GƂ�D"��۴�;�9E�iĂ ��ii�Fm��\���bn����F�RFףƧGt��ƳS�Ə��D@(�F�����<b�L��ǎÃF*�D��^Ĺ�$FY���/�r��]�����F�]2ƅX�G��Cǘ�$G���1ޙF�kG8n�E�	F�[(���1 )ǘ��G���Ħ��f��ǓW��JlFL��F	[C�����M�F\w�ī<`�d�,�(�4E�29�кD�ԚE�~F�];��L�D�>�#.�Ģ�E#$BF��p�dZĘ�?�,�^��E �f��
�.`E�=C�u���4F�pfŉP4� K@�!=F��W��j�ƅ��E��F�h"�"eF�F*İ�ŷÕE�PhEz:,Fs�����!D�3����'F�eUń_z�Ύ�F��E 2��e���\�H�Ɗ�Ŕ�e�ćV�Ŗ8�FP�]D��bFQ���D�ZC�b*L       
categories[$l#L       +                          	   
                               	         	                                                  	   
             L       categories_nodes[$l#L                      )   .   0   7L       categories_segments[$L#L                                                         )       *L       categories_sizes[$L#L                     
       
                                   L       default_left[$U#L       }                                                                                                             L       idiYL       left_children[$l#L       }               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c   e   g   i   k   m   o����   q   s   u   w   y   {��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       }O�#P�شP�U�P���Q(�:Q@�P�P��~P��1Q&p�QH�P�y>P��5QH�hP��PȣQP��P��^Q�2Q?|�Q7��Q/DQ2ƨQ��Q(��O��dP��FP>pQNtP��^P�Z�PJ�O�TO�`�PcV�Q��tP��tQ�D�QA�dP��LO@�P�ASQ9|P��P5;2P��O��NP6l~P�}WP�XPw�tOq�Oy�P͆�Of�O�`    QKVO�� P��PI�jP�P���                                                                                                                                                                                                                                                        L       parents[$l#L       }���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   9   9   :   :   ;   ;   <   <   =   =   >   >L       right_children[$l#L       }               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d   f   h   j   l   n   p����   r   t   v   x   z   |��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       }>�1'>��=��`=��>vȴ>�ƨ>oBfff?��=���A�  ='�?;d@@  D� @�  =   B�  =��BP��A�  B0  >��H      Ap     B��q@�  <�B��>;dZB�33@�  >w��>Ƨ�B�  B�  >��@�     D�@ D�@ @�  BB�R   B��q   @�ff?/�@@  D�` A`  B4z�   Ħ�D�` D�� >VB��<�`B>����M�F\w�ī<`�d�,�(�4E�29�кD�ԚE�~F�];��L�D�>�#.�Ģ�E#$BF��p�dZĘ�?�,�^��E �f��
�.`E�=C�u���4F�pfŉP4� K@�!=F��W��j�ƅ��E��F�h"�"eF�F*İ�ŷÕE�PhEz:,Fs�����!D�3����'F�eUń_z�Ύ�F��E 2��e���\�H�Ɗ�Ŕ�e�ćV�Ŗ8�FP�]D��bFQ���D�ZC�b*L       split_indices[$l#L       }         
   
         
                                                                                                                                                                                                                                                                                                                                                                                                                                      L       
split_type[$U#L       }                                                                                                                     L       sum_hessian[$d#L       }F�` FX Fh F D� CR  E�@ B@  F\ C�  CI  C
  B�  B�  E�  A�  A�  E� E�p B�  CG  C2  A�  A�  B�  B   B   @�  B�  B@  E�� AP  Ap  A  A0  C�� E` E� C+  B�  @@  B�  B�  C-  @�  A�  @�  A`  A�  Bt  B8  Ap  A�  B  @�  @�  @   B�  A@  B  AP  Cp  E�  @@  A   @�  A   @�  @�  A  @   C�� A`  D�  D7� E�� C�� C  AP  A�  B�  @   ?�  B4  B8  ?�  B�  Bh  B�  @�  ?�  A  A   @   @   A@  @   A   A  BL  A   A�  A�  A@  @@  @�  AP  B   @@  ?�  @�  @�  ?�  A�  B�  A   @   A�  Ap  @�  @�  CY  A�  D�� E�H L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       125L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       q@�3�CGH���hDiWy�1��Ľp}�o\�Dv����+�7�GD;kd�X4�Eo�%ţ����h��5D�C�G`�ǝ���a%SF��BDs:����~n�F�s�Fr�3��
qF�tƆ��OFN9zG	���G�;Dk��F��UFsX�ŉ PDzS�ǵޒF CŖ��GK��ĥÉB�@�F���"{�h#��ؾ���QG,J�ţh`�v@F�K�[�F��G6n(E/L`�vk����Ŏt��5(�Ɲ$E-W-C�����7E�OE�1�6���m���#ź�YEq�DL~g��UE�uG]��FHa�DW1
�a�&E�سC��g�
��ƒ}���l9E@�D'���j�\ŤT�C�uF���j����"�FhE�6��|FD�y�Fy�Bh�D7��Fn��Ct�3E��gF�@�EX����AEU��Ō9>ōlZ�-�EiD��y��F2�ƒ4�L       
categories[$l#L                 
                                                         
   L       categories_nodes[$l#L                                   (   -   2   :L       categories_segments[$L#L                                                         	       
                            L       categories_sizes[$L#L                                                                                           L       default_left[$U#L       q                                                                                             L       idiZL       left_children[$l#L       q               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;��������   =   ?   A������������   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c   e   g   i   k   m   o����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       qO���PuPKH|P��P�4�P@��P�P��Q��Ql^P��P[*P�yeP/�APn�HQ6��P�V�O�R�P�<Q��QV=�P��`P��P5[JP>aO�P��O��5OI�$P"        P_L�P�f�P��            N���P���Q#�bQ>.
P��-P���Q*$�O���Qt�P�u�P��P�ȿO�jP`ߣPl՜P bP��N@ܠOM��O�N�6�O�=�P2
�                                                                                                                                                                                                                L       parents[$l#L       q���                                                           	   	   
   
                                                                                                                             !   !   "   "   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <L       right_children[$l#L       q               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <��������   >   @   B������������   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d   f   h   j   l   n   p����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       q      B�     @   A�  >�$�<o>���?�{@�D�  @�  B�  =���='�B�     @@  =��   ?4��D�  D��    D��       D�� B>�FN9zG	��>��B�  >�^5FsX�ŉ PDzS�=�P=�C�   B�ffB���Bfff?Vȴ   @�  A�  @�  @�     B�  @@  =�S�>�ffD�  >fffBe33   >1'@   Ɲ$E-W-C�����7E�OE�1�6���m���#ź�YEq�DL~g��UE�uG]��FHa�DW1
�a�&E�سC��g�
��ƒ}���l9E@�D'���j�\ŤT�C�uF���j����"�FhE�6��|FD�y�Fy�Bh�D7��Fn��Ct�3E��gF�@�EX����AEU��Ō9>ōlZ�-�EiD��y��F2�ƒ4�L       split_indices[$l#L       q                      	                                              	                                         	                                  	                               
                                                                                                                                                                                                                                   L       
split_type[$U#L       q                                                                                                     L       sum_hessian[$d#L       qF�` Fx( D�� F	T Eݨ D�` B�  F	( A0  E/P E�  Dd  C�� B,  B   Ap  F� @�  @�  E)� B�  E�  A�  D_  A�  B�  Cb  Ap  A�  A�  @   ?�  A`  F, B@  @@  ?�  ?�  @�  C  E� A�  Bd  Eq@ C�  A�  A@  D� C~  A0  A  A�  B�  CQ  A�  @�  A0  A@  A�  A  A�  A0  @@  F� A�  B0  @�  ?�  @�  B  C[  D� D� A�  @�  BH  @�  D�  D�` C  C�  Ap  ?�  @�  @�  C� C+  C  B�  A   ?�  @�  @@  A`  A  B  B4  B�  B�  @�  A0  @   @   A  @   @�  @�  A  @�  @�  @@  @�  A`  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       113L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       q@�ŰD+����,D����������D2
Õ�nE_]Ɣb�D�������ɐF�'=D"�邪���AE�q��0�FMX.���F+�ƛM����$F�qm�����eOY�
�}D���C8ƕ��ǘM��!�E"7
F��E����n����ّGN������F���ĴHnF�ی�d|a�9�@�9��E�U��ע�H�Ũ��G7>ĝ��Ǔnc��LĻ�{E����+$�A���F��F����b�����,�4Ų��E���qէEiiHE�C��.=
E���į^��%�F�&D�\�ƀ�F�)F�_G����S�F97��o�ą	�GxE�6�F�k�Ʒ�F(HŪ�2E� u��5�T� E3��L�F��w2EZ G`����D��F�
'ů��FK���"�0§h��۠��<���rjX�f·Ew/gE��xC��1ã.�E�2L       
categories[$l#L                    	                                      	         L       categories_nodes[$l#L          	         #L       categories_segments[$L#L                             	       
L       categories_sizes[$L#L                                   	L       default_left[$U#L       q                                                                                                L       idi[L       left_children[$l#L       q               	                        ����            !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c   e   g   i   k   m   o��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       qO���P��_P�U*P���Q>W�Q{�BP��_P�bQ"�5Q0$�QE��Q`�Q��'    P�c�P�t(P���Q��Q�P��xQ8�Q)R_Q?q6Q
I�R#��P?jQ=��Q+�\P�?SQ2�Q7��P!��O�ȶQIbFQ��dQSYLQ��-PR/�P��QW�tQB�P��HQX�Q'�P]8�P�)�Q!��Qr|VQ�xNPT� P�0P�0QQ:4P���P�)|Qr8)P�>                                                                                                                                                                                                                                L       parents[$l#L       q���                                                           	   	   
   
                                                                                                                                   !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8L       right_children[$l#L       q               
                        ����             "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d   f   h   j   l   n   p��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       q>N�A@  ?�bND�` A   B�  ?!G�C  >��#   >_;dB�(�   F�'=>aG�?>�R   >�{@@  B`  >ۥ�>q��A`  @�  ?4z�@��>��9?�dZ>���?��D?6B�  @�  >Õ�@���   B���BI��?���B  ?��
D�  B  >�ȴ>�
=>��#?��??}D�� D�  ?�9>F��=�"�D�  @��H?�O�AP  A���F��F����b�����,�4Ų��E���qէEiiHE�C��.=
E���į^��%�F�&D�\�ƀ�F�)F�_G����S�F97��o�ą	�GxE�6�F�k�Ʒ�F(HŪ�2E� u��5�T� E3��L�F��w2EZ G`����D��F�
'ů��FK���"�0§h��۠��<���rjX�f·Ew/gE��xC��1ã.�E�2L       split_indices[$l#L       q                           
                              
         	   	               
         	                            
      
            
   
      
            	                                                                                                                                                                                                                                               L       
split_type[$U#L       q                                                                                                             L       sum_hessian[$d#L       qF�` E� F8 E�@ C�  Ex� E�0 E�p E1� CP  C�  Ep� B�  @@  E� E�� A�  D�� D�� B  C+  C<  B�  Em� B<  B�  BP  C~  E�( E�� B�  @�  A�  Dk@ C�� D  Dn  A�  A@  C  A�  B�  B�  A�  B\  EU� C�� B  A0  B�  A   A@  B   Bh  CD  D�  ER@ E�p @@  @�  B�  @�  @   Ap  @@  D  C�� C�� A�  C�  C�  D`� BX  A�  @�  A  @@  B0  B�  A�  @�  B�  ?�  Bd  A�  A�  @�  A�  A�  D�  E0 C�  Ap  A�  A�  @�  @�  A�  B,  @�  @�  @�  @�  A   B   A�  B  B�  B�  C�  D�  EO  BP  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       113L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       {A,����uCnO�	\D��E��B��TD� ��qaaE�'����Fj^��mc�}��C�R2�7�XF�.aƬ�F+�lF�X����)آF���E�v�G5��Ɛ��G��������'Di���*7��{����`���G"�F~�4��u�G��Ei�5G��F����p�|��0h�ٶKƧb"Ge�FD%���G��VF�������F>
gF��Ea�Ɣ�eǔ�eF��^ŗ�9��wD�%�E���Ĝ�����E�G��S"ET�[�v`�Ɲ�F� ~Ft�Ft���|�LA��P��F�L�=d�ŕ_��fp�N�fF/�FV9D�~�E>��G7�4��r�F.�uE�Oć�ƛJ�ú5�FgfM�5̋F�<�D�Tg��E��y�.��šWF��G�=�F ��ŝ-��>Z����F!S�ƃ��D����yg�!J�$���f�F�8C���Ų�E�c�ŬL]F�!C��fE�H�ĠBR�}D�nL       
categories[$l#L       !                                        	   
                                             
         	         L       categories_nodes[$l#L       	   	            !   -   0   2   =L       categories_segments[$L#L       	                                                                L       categories_sizes[$L#L       	                                                               L       default_left[$U#L       {                                                                                                             L       idi\L       left_children[$l#L       {               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c   e   g   i��������   k   m   o   q   s   u   w   y������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       {O���P���P:dP��$PϤ�Q�k�P	MPP�_�P�MFQ��P�aiQ�0Q�Q*��P��P?i�QC�;P݆�Q��Q�Q�
P�ijP��QUqQ��QPOO��P�t�Qw�P���P�O�P���PC�FO�,XP��xP��5P�dDP�-P��P��"Q��QP
LQ&�P�J�Q'=�P�I:P�!�Q]�QWSRY�PE�7P�TQ6�%        Pdm�P���P��P���QE��Q�MNQ=p(P�Հ                                                                                                                                                                                                                                                L       parents[$l#L       {���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   7   7   8   8   9   9   :   :   ;   ;   <   <   =   =   >   >L       right_children[$l#L       {               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d   f   h   j��������   l   n   p   r   t   v   x   z������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       {=�
=>-V=�x�B@Q�>��@�\)=8Q�B#
=B�33   B�  ?�B�  >�b   D�  =�
=?      =�\)>&�yB���D�` B�33@   @3o   >|�=D��D�  D�` D�` >�9X   =��@@  @{�@�  B�  B���D�� >��@ �9D�  @@��   >��>%   A�     ?�@��F��Ea�<���@N�R>#�
@�  =�{D��    Bx  ����E�G��S"ET�[�v`�Ɲ�F� ~Ft�Ft���|�LA��P��F�L�=d�ŕ_��fp�N�fF/�FV9D�~�E>��G7�4��r�F.�uE�Oć�ƛJ�ú5�FgfM�5̋F�<�D�Tg��E��y�.��šWF��G�=�F ��ŝ-��>Z����F!S�ƃ��D����yg�!J�$���f�F�8C���Ų�E�c�ŬL]F�!C��fE�H�ĠBR�}D�nL       split_indices[$l#L       {      
         
                                                                                            	                                       	             	   
                                                                                                                                                                                                                                                                                 L       
split_type[$U#L       {                                                                                                                  L       sum_hessian[$d#L       {F�` E� Fj� C�� D�` C�  Fe B�  C.  C�� D�@ Cl  B�  C�� F], B�  B<  C  B  C*  C  D�� B  C6  BX  B�  @@  Bx  Cހ F, E�  B<  A�  A@  B  A�  B�  A�  A@  B�  B�  A�  C   D�@ B,  A@  A�  C  A�  A�  B  B�  A�  @   ?�  BP  A   B�  C�� C+  E�  C� E� A�  A�  A�  @�  A   @�  @�  A�  A  A   Bt  Bt  A`  A  A0  ?�  B4  A�  B�  A�  A�  @   B�  A0  C`  D�@ A�  A�  @   A   A`  A0  A�  C  @@  A�  AP  @�  A�  A   B�  @�  A�  @�  A�  B  @�  @@  A�  BT  C�  B�  B  C
  A   E�� Cg  Cv  E� C�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       123L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       oA<�����C#ř�hE�&�Bi�TE���zƎҞEZ|"G>��Ŕ?CqǟEY�G� ����E�VZ��FB��TF�FN{F�1-G�Q�D�K@�I%�Y�|C���F��d�%�gF�4 G/��ſ8��Ax�F�����Ƃ5��t+��{;�G�]����{F�T�G#��C�ĺ�
��G	|�GGE��tE���ƒ
zD1ϣ��c}ƚ ŜH#GW�C��F�SG�J�EL����]�Sk FI0o�A^��� DK'�Fr�ňIƇ�YE>������@����)V�D�d-���F�n��6BEF�R�g�+F�2g�y��F�%�F����%�DG����F]�D�����e�E%�F���&�E�˪�9��Ű&��ھ��O�oD��F�e�E c�_7�D;�E��ƕ�4EЇ�G9��ɬ�F�E�D'1��$�dďX�ő>ML       
categories[$l#L       &                                                       	   
                                           	   
               L       categories_nodes[$l#L       	   #   &   (   *   +   ,   2   5   ;L       categories_segments[$L#L       	                                           	                     %L       categories_sizes[$L#L       	                                                               L       default_left[$U#L       o                                                                                                   L       idi]L       left_children[$l#L       o               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;����   =����   ?   A   C   E   G   I   K   M   O   Q   S   U��������   W   Y   [   ]����   _   a   c   e   g   i   k   m������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       oO�VLP�bPP&�?P�pJQ$�PO}�Q^hP��GQA�Q	��Q�P��:P%.4Q�Q+pR
��Q,�=Q�~QA�^Q	&QC5Pa��O
�@P���Q�PP�,�P�,�QrfQ01O���    P��    Q�>�PW]<P���Q7�ZP�^P��tP��P��QqbQ���M�|�O��l        QaQ2��P��QM��    P��P(��P �P�LP�u�QQ�u�K�k�                                                                                                                                                                                                            L       parents[$l#L       o���                                                           	   	   
   
                                                                                                                           !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   /   /   0   0   1   1   2   2   4   4   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;L       right_children[$l#L       o               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <����   >����   @   B   D   F   H   J   L   N   P   R   T   V��������   X   Z   \   ^����   `   b   d   f   h   j   l   n������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       o=49XD�  B�  >���A�  ?=p�>   >R�D�  >��^>���>�JD�  =e`BB8��>O�;?u?�dZ?o�;@�p�B4z�>oB���?(��BH>��9D�@ >P�`B��{@   G/��@����Ax�@��>���   D�` @@     @�     B�
         GGE��t>\)D�` >�   ƚ @      B��D�  @@  B�  D�@    FI0o�A^��� DK'�Fr�ňIƇ�YE>������@����)V�D�d-���F�n��6BEF�R�g�+F�2g�y��F�%�F����%�DG����F]�D�����e�E%�F���&�E�˪�9��Ű&��ھ��O�oD��F�e�E c�_7�D;�E��ƕ�4EЇ�G9��ɬ�F�E�D'1��$�dďX�ő>ML       split_indices[$l#L       o                                    	               
               
            
                                                                                                                                                                                                                                                                                                                            L       
split_type[$U#L       o                                                                                                      L       sum_hessian[$d#L       oF�` D�  F{@ D[@ Cs  Fw` Cx  D5  C  C]  A�  D� FnH Cn  A   C�  C�  B�  A�  B�  C  A�  @�  C�� Cs  BX  Fmp B(  CD  @�  @�  C�� @�  C�� B  B�  A�  A�  A   B|  A�  B,  B�  @@  AP  @�  ?�  C�� BX  B�  B�  @�  B<  @�  Fm\ B  @�  C&  A�  @@  @@  C�  B|  C�  B  A�  A0  A�  B�  A�  @�  A   A0  @   A   B4  A�  A   A  A   B  @�  B�  @   ?�  A  @�  A�  C~  @�  BH  B  B�  B�  A   A  B  @   @@  FO� D�` B   @@  @@  @�  C  A@  A�  @�  ?�  @   L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       111L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       }A�ZC�����C�՝Ţ��c��F\��B�E�O�<��F���FS��Ǧ���4G'�ţ1�C��GF��(�n$�ƝI�E�}�F+��Gg��F�X��N�8�FP�Aǡ#'E}�EƨsG�+m�N6��lZC:8E���F���
~����ǦN��X*mǔSG����G �;E�,Fi��GژdE��G$X��SX�;ADӷA�:#MFѝ3�']�Ţ؀�#dG	2'�瞲G�7m�8iFW	G�rC�?�� �'D����B�6r�EwoD1�7F��	E;��FN�WE�.A�"�ŵ�dE�r�EN��Be1E������g��~�E��fF��EE/�ŋy�F���EJvF��Ķ=�FIFܝb��BG$�����R�iE��G5�sF#�%D�=S�#Ed��4�t�
Ħ�F#��D�mŚ��FK
;��\�ƵlzŞ�2E.m���Fq��^����ĂŚ�NG>wD�^�E�z�&�{Fɖ��;�~GH��)�L       
categories[$l#L       4      
                	   
                                                          	                               	   
                                           L       categories_nodes[$l#L                          &   '   )   .   4   ;L       categories_segments[$L#L                                                                       )       *       3L       categories_sizes[$L#L                                                                             	       L       default_left[$U#L       }                                                                                                           L       idi^L       left_children[$l#L       }               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c   e   g   i   k   m   o����   q   s   u   w   y   {��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       }O���P0GwP�̝P�rsQ�ݰQ2^Q<&�P>�Q�#JQ9YyQ �#Q�HQ
eoQ+��QTw�P�b�PH:Q��Q���Q���Q�6P6c,Q'�PQA%�O�P�bVQv�CP��QJ�\Q�QQ�e�P���Pթ�P���QH�*Q3#$P��Q|*Q��Q=ЎP��P��$Q�O��P01RQ
�PֽlP�MfQ�OUӴO.��QQ,?>Q�9PO�N��L    Q�@P���PN{�Pk^�P:�GQ~��                                                                                                                                                                                                                                                        L       parents[$l#L       }���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   9   9   :   :   ;   ;   <   <   =   =   >   >L       right_children[$l#L       }               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d   f   h   j   l   n   p����   r   t   v   x   z   |��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       }A   A@  B�  @�  >���D�� @��?
=q?�5?>�G�By33   D�` D�� D�� >�ffB�     @�  >�bNB$ff>���?X��B9��B{?-�h>���      @�  @�ffB�
=   B�  @�  B:ffBL  ?\�      B0     B���B  @�>1'   >fff=ix�>�P=L��D�@    >��/>��7D�� �#d>vȴA     A@  >.{@JC�?�� �'D����B�6r�EwoD1�7F��	E;��FN�WE�.A�"�ŵ�dE�r�EN��Be1E������g��~�E��fF��EE/�ŋy�F���EJvF��Ķ=�FIFܝb��BG$�����R�iE��G5�sF#�%D�=S�#Ed��4�t�
Ħ�F#��D�mŚ��FK
;��\�ƵlzŞ�2E.m���Fq��^����ĂŚ�NG>wD�^�E�z�&�{Fɖ��;�~GH��)�L       split_indices[$l#L       }                              	                                	         
                                               
                           	                            	                                                                                                                                                                                                                                                                                 L       
split_type[$U#L       }                                                                                                                  L       sum_hessian[$d#L       }F�` Fz� D�� Ft< Cɀ D�� B�  Fn0 C�� C�� B�  C8  D[  B`  BH  Cـ Fgd Co  C  Cd  B�  Bl  A�  C  A�  DE� B�  @�  BH  A�  A�  C�  C  Fd� C(  C2  Bt  C  A@  CN  A�  B  Bx  A   BD  A0  A   B�  BX  @�  A�  CE  D� B�  A�  @@  @@  A�  A�  @�  A�  A0  A0  C�  A�  B`  B�  Fd� A@  C  Ap  B�  B�  A�  B  B�  B$  @�  @�  B   C&  A�  @   A�  A�  Bl  @@  @�  @�  B  A@  @@  A   @�  ?�  Bl  B8  @   BP  @�  @@  @   A�  C'  A�  C   C�  B8  A�  @�  A   @   ?�  A�  @�  @@  A�  @@  @   A0  A@  ?�  A   A   @@  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       125L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       wAU0�CV�&ı����/E��xűG�EM��}؎D5�zFt0>�]��� ���¥[D��dF����'�O	��Q�D�aPE�x�G2?F��_��(�G�F� �ƆbǞ+�D�8�@��k�VG]�LF<��,�b�����7�$E>9�ŏ[3Gh��D��JG�93E���ƫ��GK��E�:Gw��e{�ņ&4��u~ưQ�E|�C���
cFƌ��D@�F�����������fn�MCG�>�S&�F�Ź:ą� B��x�Y�E��AF�Îƙ'��iE����&�C�mF�qAEz]�D�G�C1UGX��Ĝ�E��m�8��FK���x�F���DeT��>ոFG{�F��C����(��V�=C��*�ޝC�3��<{h�6��Eq�M��E��/ƍ��Ů��L��3iE\d�ƾ�D�x[Ģ%�Fh'N�!�.�c��F���u3��.n�F:�ų�ME�4G ���	3~E�:�L       
categories[$l#L       )                         	   
                               	   
                                           	   
                   L       categories_nodes[$l#L                    %   '   8L       categories_segments[$L#L                      
                     %       &L       categories_sizes[$L#L              
                                   L       default_left[$U#L       w                                                                                                        L       idi_L       left_children[$l#L       w               	                                    !   #   %   '   )   +   -   /����   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c   e   g   i   k   m   o   q����   s   u����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       wO���P��P�d�P!9#QG`�QV�;Pݐ�QK5Pr�yQgJ�P۵/Q*��QS�vQ,�GQ��P{~�Q5��P�Q�UQ�"Q��^P�XFQ$�Q(O    Q.QZqP��<Q8��Q��QIeZQḍP��P�d�Q�>9Q.ÂP�8aQ-?ZP�pTP��P�P�Q UQ�t$P}nQP�P��P���Q8�Qe��Q&P�7TO�)@P���P���Qp�{P�?OO��0O?W�    Q��O��A                                                                                                                                                                                                                                        L       parents[$l#L       w���                                                           	   	   
   
                                                                                                                                   !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   ;   ;   <   <L       right_children[$l#L       w               
                                     "   $   &   (   *   ,   .   0����   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d   f   h   j   l   n   p   r����   t   v����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       wD�� D�` ?H��>_;d   ?*~�B�  >Xb>��B~=q? �?�|�B��=B�(�>7K�   B�� =��? A�=u?S�F@Dz�?Fff@�ffF� �@S�
@�  @�  ?;"�@���B�ff@�     >�ȴD�� =��w>��
   ?�z�   BDff>/�?���@�  ?u@@  @�  ?>�R@I�?/�>��^?�z�?y��@@  >���@@     >o�MC>�ȴB�  F�Ź:ą� B��x�Y�E��AF�Îƙ'��iE����&�C�mF�qAEz]�D�G�C1UGX��Ĝ�E��m�8��FK���x�F���DeT��>ոFG{�F��C����(��V�=C��*�ޝC�3��<{h�6��Eq�M��E��/ƍ��Ů��L��3iE\d�ƾ�D�x[Ģ%�Fh'N�!�.�c��F���u3��.n�F:�ų�ME�4G ���	3~E�:�L       split_indices[$l#L       w         
          
                  	                         
                            	                                        	   
      
                                                                                                                                                                                                                                                                                          L       
split_type[$U#L       w                                                                                                                 L       sum_hessian[$d#L       wF�` Fk� E0 Fb� D@ Dq@ D�� E�� F 8 C�  C�� DP  C  D�� B  E�h C�� D�� E�� CM  B�  B0  Co  DN� @�  B�  Ap  D�� A�  A  A�  B�  E�  Ci  B  D� D�� A�  E�X @   CK  A�  B�  B   A@  Ap  C`  D4� B�  B<  B�  @�  A   D~� B�  A0  @�  @�  @@  A�  A   B�  B  D�  E�  CQ  A�  @�  B   C�  B�  D)@ C�  A  A0  D�  E�� ?�  ?�  B�  B�  @�  AP  B8  A�  A�  @�  A   @�  @�  A   C8  B   D-� A�  B�  B  A�  A�  A�  BL  ?�  @�  @�  @   C�  D@ B  B  @�  @�  @@  @@  ?�  @�  @�  Ap  @�  @�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       119L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       w@���B��1�$ՠ� )�D�2gEA<*���CP՞�Ay�ŪZ*Eb�G
7�kZ��N��Fvx�ԁE�}n��
>�"�E���g`�Ŭ�E���GJ�/�ƕg��D�jN�n���Gm�(E�z���Ʊg5FFΨ��P�E $�1D�ƫ�m�Y��ŷ�QF�s��2İ��ƹ�O�G�E�����Gu����r�Ę� Ƨ����rF���T0s�T��F�+g��u��K?�F�ΒE���FV����xC71m�A��aS�D�m��O+�E�Ҭ�H}rF�;�BS'Eqp0E`4�ŵ�HD���E�8Ť�f��Ƨ�AF��EO�aD�	��'���!� �<f(�*QE����7f�Ej�
��%_F�0?��lE+�ƽ�
D7
gF����9VS�2g�AL�7�j��ɱF? �7�D���E�@�Še�E�Fr]CE*�#�ٿ�Ƙ��Ĝ��� ��F4.E��m�2�L       
categories[$l#L       9               	               	                                                    	   
                                        	   
                                                     L       categories_nodes[$l#L             	   
                  %   &   '   -   /   >L       categories_segments[$L#L                                                                -       /       0       5       6       7       8L       categories_sizes[$L#L                                                                                                         L       default_left[$U#L       w                                                                                              L       idi`L       left_children[$l#L       w               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c��������   e   g   i   k   m   o   q��������   s   u��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       wO�k�Oً�P�z�P`/~Q�wQ&��P̣�P���Pݻ�QW��Q#IMQ�-P���P��$PXs-P���Q8�}P�BP�6�P�KQ�VQt>Q��P�{4M�)�Ox�P��P��\P`~pN���O�7BP�;�P�$fQa��Q�P�]�Q�|P�B(Q�sP�P���P��EQ�P�~QoWQ���P�OO��P�tM]%�        N�̀Q4	�P?LP�]�P�mOW�PR.�        O�`�Oruy                                                                                                                                                                                                                                L       parents[$l#L       w���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   4   4   5   5   6   6   7   7   8   8   9   9   :   :   =   =   >   >L       right_children[$l#L       w               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d��������   f   h   j   l   n   p   r��������   t   v��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       w?��@�   ?��D�� ?}�-D�  ?-B���      A$��>�  @�Q�   ?�n�?,I�   D�� >�
=@@  @��
   >��A)G�>H�9?��?�t�B0�\      @��@@  @�Ap  Bk��B"           >BF��>_;d?A%>�ȴ   @��   @�  D�� Ę� Ƨ�@�  B`\)@�  >oB���@��D�� F�ΒE���?�;d   C71m�A��aS�D�m��O+�E�Ҭ�H}rF�;�BS'Eqp0E`4�ŵ�HD���E�8Ť�f��Ƨ�AF��EO�aD�	��'���!� �<f(�*QE����7f�Ej�
��%_F�0?��lE+�ƽ�
D7
gF����9VS�2g�AL�7�j��ɱF? �7�D���E�@�Še�E�Fr]CE*�#�ٿ�Ƙ��Ĝ��� ��F4.E��m�2�L       split_indices[$l#L       w   	                      	                            	                       
                                                                	                                                          	                                                                                                                                                                                                                                   L       
split_type[$U#L       w                                                                                                         L       sum_hessian[$d#L       wF�` F�� D9  FY  E � C�  C�  F@� D�� D
� D�@ B  C�  C�  B  F2 Dk@ D�� Cˀ C}  C�� C�  D�@ A�  A   A�  C�� C~  B  @�  A�  F1� B  C̀ D  Dh  CW  C  C  B�  C   C
  C#  B�  C�  B@  D�@ @@  A�  @�  ?�  @   A�  B�  C�� Ca  A�  A@  A�  @@  @   A�  @�  F� E� A�  A�  CA  CX  D@ @@  DF  C  B\  C   A�  B�  C  B�  B�  @�  A`  B�  B�  A�  B�  B�  B�  A�  C7  C  A�  A�  D$� D`  ?�  @   A�  @�  @�  @   A`  @@  B  B0  C  C  A�  CI  A�  @�  @�  @�  A�  @�  AP  AP  ?�  @�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       119L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       @�ðC�wO�\VD��FĜ(��¶�DF�5DNC�FY�;D����\إE��������E�tD�͎�˗@Ƌ
Fޮ��w_nFZd���ġ��F����f���u�ƝyE~����Fl��
Į�E�z�(����>G	���G(�E�ao��Z^D�a#F�h$�!�ƛ��EXG�Et�����DM�Gm��-FeF�t��oRG��#�|ED*�*���E�aE���š~�G��FG����E�|�D���Ďk?��DHiGF;@ĵ�0Fܴ�$E��˝�Fη�ų���>>E�u`F�:��9��E�c*�D�qD�ޅD����JE��F�ƶa�D�%l���E "�CށvG!�9C�H�F)��7�]ņ��Ff���m"�F?�F�M_���C���SFg�l� ��~;�5���S��F��F��U�2*�F6x��^8ï�.��O�Eq��� ��Ć�EU�S�!�Ca��G�8E���E�՗��V�#E�cC�E�pŇ�	L       
categories[$l#L                         	   
                               	                L       categories_nodes[$l#L                "   )L       categories_segments[$L#L                      	              L       categories_sizes[$L#L              	                     L       default_left[$U#L                                                                                                                     L       idiaL       left_children[$l#L                      	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c   e   g   i   k   m   o   q   s   u   w   y   {   }����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       O��P�h�Q'sNQ"b�P�G�Q��QwPs�Q�w�Q@�P�O�Q.��P�tP�w�Q�UP��P�ՊQ��'Qo8QXmQ8,NQ�5�Q#��P���Pp�2Q��NQW�>Q3_Q,M6Q0*�P���P�]P���P�ftP��QQ�#�Q9��Q���P�k�Q(�Q� QD�QP�Qa$XQ���Q\��P�$�P�-�P�<PP�kPsѷP��P���P�6�Q�(�PЇ�QDD(Q��P���P��Q2��P�l�QP��                                                                                                                                                                                                                                                                L       parents[$l#L       ���                                                           	   	   
   
                                                                                                                                         !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <   =   =   >   >L       right_children[$l#L                      
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d   f   h   j   l   n   p   r   t   v   x   z   |   ~����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       @�  D�� @�  D�` ?�33>�P@bN@7�w?	7LA��>�
=   B�     @�  >1&�B�  >k�@��HD�  >���@,�@.v�BS�H>��TB�  D�` =�x�>O�@I�>;dZB0  A�R=�j   Bq33B���@o=�G�>��T@��   >��#@�  A0  @'�?*=q>��>�-B[z�D�� B�G�@"�\>L��>�S�Be33>��D�� @�=q@�  ?	�^?��>�A�D���Ďk?��DHiGF;@ĵ�0Fܴ�$E��˝�Fη�ų���>>E�u`F�:��9��E�c*�D�qD�ޅD����JE��F�ƶa�D�%l���E "�CށvG!�9C�H�F)��7�]ņ��Ff���m"�F?�F�M_���C���SFg�l� ��~;�5���S��F��F��U�2*�F6x��^8ï�.��O�Eq��� ��Ć�EU�S�!�Ca��G�8E���E�՗��V�#E�cC�E�pŇ�	L       split_indices[$l#L                         	      
   
                       	      	         	                                                                  
                                                      	                                                                                                                                                                                                                                                                      L       
split_type[$U#L                                                                                                                                  L       sum_hessian[$d#L       F�` F>� E�� E�p E�� D�` EnP E�H C�� D�� E� Cm  Do� EJ� D� E�0 C�� B�  C3  D�  Ce  D  DӀ B�  C  D@� C;  De� E� C�  Ch  E� E�p Cw  B0  A�  Bh  B�  B�  B�  D�  C   B�  C�  C�  DN� DX@ B0  Bp  B�  A0  D>� A  B�  B�  CJ  D3  D,  D�  A0  C�� B�  C  D&@ D�� CD  E�P A0  Cl  @�  B  A@  A@  B   A�  B�  B<  AP  B\  B`  B   D�� C�� B�  A�  A   B�  C�� Bt  C�� @@  DA� BP  D@ C�  A  B  B`  @�  B�  B<  A   @@  D6� A�  @   @�  @@  B�  B  B4  C  B�  D  C4  C�� C�� D�  D@ @�  @�  Cc  B�  B�  A�  B�  B�  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       127L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       uAܢ�p"E%|W��,C�
^F��ħE��x�Eoc,B��E����p�FD^$�6�"E���n��(WNF�	uC�:i�-i�F�k��T�HFF��EV���+	�F�`�E��RƊ��E��G/�GDؼ�Ğ��Ƴ��Ʀ�>D��DGR	 Ƈw.F
QO�	ɊÈ��E� �G�9�E�:��	A�F�tF�j��j��Ɛ$�F���ǽH�C�FÅkGh��kgF�d��#�D�C4mG<|���wF	��Ńw��IIŁ�E����9���ٖ�F�7bF"�8Ĩ6 G`eyF:!VDE���V�����%E�G�D���$B9��ă�E[������FϘC��4E�±�N��i$D�h�F����#�F.��E��E3�,��C���2�Ɵ��5��F���Y��E�O�I��F��7D����5��F�n�F�V!E�8��k��L[dƹ��ű�Fێł�cE�۠�Gj�"`�Ţ}1L       
categories[$l#L       6                      
                                                 	   
                                     
                               	   
                        L       categories_nodes[$l#L       	                        #   -L       categories_segments[$L#L       	                                    "       %       3       4       5L       categories_sizes[$L#L       	                                                               L       default_left[$U#L       u                                                                                                    L       idibL       left_children[$l#L       u               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9����   ;   =   ?   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c   e����   g   i   k   m����   o   q   s��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       uO�FlPY7�P�ɪPͨ.P���Q	ݎP�j�P�ZDQ$H:P��Q��P�%�Q-r�P�H�Q"�P���Qce�Q�7�QqP��!P�l�Q��Qe�P��9Q��Q��fP�aCP�HQ:�[    P�6�P�@�Q�Q�:Q"�Q���Pw��P�
@QMnP�>�Q��P7�P�SP�=�P�u�QV�2O�YbP5c�P�`P�P	�Q��`    P�~]P/��O��vP��@    Pm��P��4PC4                                                                                                                                                                                                                                L       parents[$l#L       u���                                                           	   	   
   
                                                                                                                                   !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   5   5   6   6   7   7   8   8   :   :   ;   ;   <   <L       right_children[$l#L       u               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :����   <   >   @   B   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d   f����   h   j   l   n����   p   r   t��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       u?WK�@�     A0  ?�P>�S�?I��      ?S��=�;d>A�7?�n�@Ĝ>� �A   @4�?;"�D�� ?I�>��9D�     >���>D��A33@�m      G/�G   ?:�B:ffA0  >�=q   Bs��?�E�Btp�>��>��@�  D�` @�  B      D�` @�  B8��@@  D�  ?�~�Gh�@�  @&B��{@@  G<|@:�\?� �D�� �IIŁ�E����9���ٖ�F�7bF"�8Ĩ6 G`eyF:!VDE���V�����%E�G�D���$B9��ă�E[������FϘC��4E�±�N��i$D�h�F����#�F.��E��E3�,��C���2�Ɵ��5��F���Y��E�O�I��F��7D����5��F�n�F�V!E�8��k��L[dƹ��ű�Fێł�cE�۠�Gj�"`�Ţ}1L       split_indices[$l#L       u                   
                          
   
         	                            
                           	                                                                          
                                                                                                                                                                                                                                      L       
split_type[$U#L       u                                                                                                            L       sum_hessian[$d#L       uF�` F}  D|  E'p FS$ C�  D� EP D� FL� Cǀ BX  C�  C!  C�� D�� C�  B�  C�� FLH B   B�  C�  B  A�  B�  Cq  B�  B$  ?�  C�  D�@ Bt  Cw  CO  B4  A�  C�  Co  FD� C�� A   A�  B  B  C�  B0  A�  A`  @�  A`  B�  @   C)  B�  B�  A�  ?�  B   CL  Ct  D�` B�  A�  B(  Cr  @�  B  C.  @@  B(  A�  A0  C  B�  C   B�  F-� D�  C�� C$  A   @   A�  A`  A�  A   @�  A�  B�  C=  A   B  A�  @@  @�  @�  @�  @@  A  @�  B   B�  C'  @   @@  B�  B�  @�  A   A0  A0  A�  B�  B�  C;  Bd  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       117L       size_leaf_vectorSL       1}}{L       base_weights[$d#L       }A��7�i�RC��DYW��2B�F9SC1��Ŗ�dEV�[�`E�mLF��
Ġ�OáDCE(�]DLy>�#7bFU�Du��E�pŌ��F��C�#�8F�m�D�fOF�ŎhDBs��6�+E���Ņ�xDܶhƞ�(�[�Ft�4F_�Ŝ�F4��C�qtD�DGc'ĂFx��W���oGF�\s�^^�G� �F�#!G��Ǌ+qE顜E矴G]�yD�B���!�C���F�T'D7�����F	I�C�6Yƛ��D0�×s5F5�Ć�o��RĽ+<F+�n�)��E����5Xfƥ��E����ĭ�XD��E1���[~�_��G�3�e��E�<��_ͭ�p�Cű�MF0�zE��F8�������M/�F잿E�oA�\�kF
\G�E�Ч�5�4ƽߑō�yEũ���"E�KFҐ�E�|2E���o�x�;W�E�CJ��5E(;�FPHD�D�� �����'�`�3F��D�PE4� ��b���JE6���P�E��ZL       
categories[$l#L       R                                             
                      
                               
                                               	   
                                         	   
                                  	                               L       categories_nodes[$l#L                               .   1   4   9   :   >L       categories_segments[$L#L                                                  "       #       $       2       3       @       J       QL       categories_sizes[$L#L                            
              
                                          
              L       default_left[$U#L       }                                                                                                            L       idicL       left_children[$l#L       }               	                                    !   #   %   '   )   +   -   /   1   3   5   7   9   ;   =   ?����   A   C   E   G   I   K   M   O   Q   S   U   W   Y   [   ]   _   a   c   e   g   i   k   m   o   q   s   u   w   y   {��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       loss_changes[$d#L       }Oѥ�P�c�P�6�P�ˢP|��P���PY>P��PP���P��KQ��Q({PK�PPͅ'P�f�P��PP�?YP�D�PA��P�/QP���Py�lPź�Q��P��2P]P{��Q@YHQHpP���Q��P�5�    Q!wPl$�P��P��zP��PT�hP��Qw��Q��P���P P��vPv��N��`P�d�P.�O1aXP��7O9�O�)@P��aPY��Q(zQ�QQN��P鼴Q2G�Q$P�t�P�է                                                                                                                                                                                                                                                        L       parents[$l#L       }���                                                           	   	   
   
                                                                                                                                 !   !   "   "   #   #   $   $   %   %   &   &   '   '   (   (   )   )   *   *   +   +   ,   ,   -   -   .   .   /   /   0   0   1   1   2   2   3   3   4   4   5   5   6   6   7   7   8   8   9   9   :   :   ;   ;   <   <   =   =   >   >L       right_children[$l#L       }               
                                     "   $   &   (   *   ,   .   0   2   4   6   8   :   <   >   @����   B   D   F   H   J   L   N   P   R   T   V   X   Z   \   ^   `   b   d   f   h   j   l   n   p   r   t   v   x   z   |��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L       split_conditions[$d#L       }B5\)   B8��   @a%   ?�@qG�>���=�9X?D�@�z�>�>��H   C  D��    =D��?�;Bff@@  @@  ?-V@��D��    >�9X>��+   @@  B2  ƞ�(D�� ?�&�A�R?ߝ�@@  @z�>`A�D�@ B  >�$�@@  >���@�     =��`@�     >�\)>�(�   ?���>ۥ�>�!>�
=      @@  @���@��   ×s5F5�Ć�o��RĽ+<F+�n�)��E����5Xfƥ��E����ĭ�XD��E1���[~�_��G�3�e��E�<��_ͭ�p�Cű�MF0�zE��F8�������M/�F잿E�oA�\�kF
\G�E�Ч�5�4ƽߑō�yEũ���"E�KFҐ�E�|2E���o�x�;W�E�CJ��5E(;�FPHD�D�� �����'�`�3F��D�PE4� ��b���JE6���P�E��ZL       split_indices[$l#L       }                             
            	                       	                                              
                        	      	          
         	          
         	                 
                                                                                                                                                                                                                                                           L       
split_type[$U#L       }                                                                                                                L       sum_hessian[$d#L       }F�` E�� F9| E+� E!p C�  F4T D@ EP E0 C$  C5  C  Fx D�� C�  C�� C�� D�� C�  EP B�  B�  B�  B�  Ap  C  Eӈ E2� D�  C�  C�� @@  C�  B  C�� B�  B�  D�@ C~  A�  Du  D�  A�  B�  B�  @   B�  A   @�  B�  A   @�  B�  A�  E�P C'  D�� D�� D@@ D.  B�  C�� C�� A�  C  B�  A�  A�  B$  Cl  B�  @@  BP  B`  Cـ D�� C$  B�  A   @�  D]  B�  D@ D  A`  @@  A�  B4  B`  A`  ?�  ?�  @�  B�  @�  @   ?�  @�  A�  B4  @�  @�  @   @@  B\  BH  A�  A  E�H B  B�  B(  D�� D� C�  D;� B�  D.  C�� CՀ B�  A�  C�  B  L       
tree_param{L       num_deletedSL       0L       num_featureSL       24L       	num_nodesSL       125L       size_leaf_vectorSL       1}}}L       nameSL       gbtree}L       learner_model_param{L       
base_scoreSL       8.2300875E5L       boost_from_averageSL       1L       	num_classSL       0L       num_featureSL       24L       
num_targetSL       1}L       	objective{L       nameSL       reg:squarederrorL       reg_loss_param{L       scale_pos_weightSL       1}}}L       version[#L       ii i}}�
       ���R�sbub.